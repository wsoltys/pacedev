-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_SND_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_SND_1 is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"5E",x"23",x"56",x"D5",x"C9",x"15",x"08",x"2F", -- 0x0000
    x"08",x"45",x"08",x"62",x"08",x"62",x"08",x"62", -- 0x0008
    x"08",x"62",x"08",x"62",x"08",x"DD",x"6E",x"02", -- 0x0010
    x"DD",x"66",x"03",x"4E",x"CB",x"21",x"06",x"00", -- 0x0018
    x"21",x"B3",x"08",x"09",x"5E",x"23",x"56",x"DD", -- 0x0020
    x"73",x"04",x"DD",x"72",x"05",x"18",x"23",x"DD", -- 0x0028
    x"6E",x"02",x"DD",x"66",x"03",x"4E",x"06",x"00", -- 0x0030
    x"21",x"4B",x"09",x"09",x"7E",x"32",x"A2",x"42", -- 0x0038
    x"DD",x"77",x"01",x"18",x"0D",x"DD",x"6E",x"02", -- 0x0040
    x"DD",x"66",x"03",x"7E",x"DD",x"77",x"06",x"DD", -- 0x0048
    x"77",x"07",x"DD",x"6E",x"02",x"DD",x"66",x"03", -- 0x0050
    x"23",x"DD",x"75",x"02",x"DD",x"74",x"03",x"C3", -- 0x0058
    x"D9",x"07",x"06",x"00",x"DF",x"DD",x"36",x"00", -- 0x0060
    x"FF",x"C9",x"CD",x"72",x"08",x"06",x"00",x"DF", -- 0x0068
    x"18",x"33",x"78",x"E6",x"E0",x"07",x"07",x"07", -- 0x0070
    x"47",x"3E",x"01",x"10",x"04",x"DD",x"77",x"00", -- 0x0078
    x"C9",x"07",x"18",x"F7",x"C5",x"CD",x"72",x"08", -- 0x0080
    x"C1",x"78",x"E6",x"1F",x"3D",x"07",x"4F",x"06", -- 0x0088
    x"00",x"DD",x"6E",x"04",x"DD",x"66",x"05",x"09", -- 0x0090
    x"5E",x"23",x"56",x"EB",x"EF",x"DD",x"46",x"06", -- 0x0098
    x"78",x"DD",x"77",x"07",x"DF",x"DD",x"6E",x"02", -- 0x00A0
    x"DD",x"66",x"03",x"23",x"DD",x"75",x"02",x"DD", -- 0x00A8
    x"74",x"03",x"C9",x"D3",x"08",x"D7",x"08",x"DB", -- 0x00B0
    x"08",x"DF",x"08",x"E3",x"08",x"E7",x"08",x"EB", -- 0x00B8
    x"08",x"EF",x"08",x"F3",x"08",x"F7",x"08",x"FB", -- 0x00C0
    x"08",x"FF",x"08",x"03",x"09",x"07",x"09",x"0B", -- 0x00C8
    x"09",x"0F",x"09",x"6B",x"08",x"F2",x"07",x"80", -- 0x00D0
    x"07",x"14",x"07",x"AE",x"06",x"4E",x"06",x"F3", -- 0x00D8
    x"05",x"9E",x"05",x"4E",x"05",x"01",x"05",x"B9", -- 0x00E0
    x"04",x"76",x"04",x"36",x"04",x"F9",x"03",x"C0", -- 0x00E8
    x"03",x"8A",x"03",x"57",x"03",x"27",x"03",x"FA", -- 0x00F0
    x"02",x"CF",x"02",x"A7",x"02",x"81",x"02",x"5D", -- 0x00F8
    x"02",x"3B",x"02",x"1B",x"02",x"FD",x"01",x"E0", -- 0x0100
    x"01",x"C5",x"01",x"AC",x"01",x"94",x"01",x"7D", -- 0x0108
    x"01",x"68",x"01",x"53",x"01",x"40",x"01",x"2E", -- 0x0110
    x"01",x"1D",x"01",x"0D",x"01",x"FE",x"00",x"F0", -- 0x0118
    x"00",x"E3",x"00",x"D6",x"00",x"CA",x"00",x"BE", -- 0x0120
    x"00",x"B4",x"00",x"AA",x"00",x"A0",x"00",x"97", -- 0x0128
    x"00",x"8F",x"00",x"87",x"00",x"7F",x"00",x"78", -- 0x0130
    x"00",x"71",x"00",x"6B",x"00",x"65",x"00",x"5F", -- 0x0138
    x"00",x"5A",x"00",x"55",x"00",x"50",x"00",x"4C", -- 0x0140
    x"00",x"47",x"00",x"04",x"08",x"34",x"2C",x"25", -- 0x0148
    x"21",x"1D",x"1A",x"18",x"16",x"14",x"13",x"11", -- 0x0150
    x"10",x"0F",x"0A",x"21",x"A5",x"42",x"7E",x"A7", -- 0x0158
    x"C0",x"21",x"93",x"09",x"11",x"80",x"42",x"01", -- 0x0160
    x"18",x"00",x"ED",x"B0",x"3A",x"A3",x"42",x"87", -- 0x0168
    x"4F",x"87",x"81",x"4F",x"06",x"00",x"21",x"AB", -- 0x0170
    x"09",x"09",x"11",x"82",x"42",x"CD",x"89",x"09", -- 0x0178
    x"11",x"8A",x"42",x"CD",x"89",x"09",x"11",x"92", -- 0x0180
    x"42",x"7E",x"12",x"CD",x"90",x"09",x"7E",x"12", -- 0x0188
    x"23",x"13",x"C9",x"01",x"01",x"00",x"00",x"00", -- 0x0190
    x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00", -- 0x01A0
    x"00",x"00",x"00",x"47",x"0A",x"6A",x"0A",x"8D", -- 0x01A8
    x"0A",x"CE",x"0A",x"E7",x"0A",x"3A",x"0B",x"FB", -- 0x01B0
    x"0A",x"19",x"0B",x"3A",x"0B",x"15",x"0C",x"3A", -- 0x01B8
    x"0B",x"3A",x"0B",x"00",x"00",x"00",x"00",x"00", -- 0x01C0
    x"00",x"B5",x"0B",x"E6",x"0B",x"3A",x"0B",x"2A", -- 0x01C8
    x"0C",x"55",x"0C",x"3A",x"0B",x"7E",x"0C",x"BA", -- 0x01D0
    x"0C",x"3A",x"0B",x"EE",x"0C",x"1A",x"0D",x"3A", -- 0x01D8
    x"0B",x"43",x"0D",x"7B",x"0D",x"3A",x"0B",x"9F", -- 0x01E0
    x"0D",x"D2",x"0D",x"3A",x"0B",x"03",x"0E",x"5C", -- 0x01E8
    x"0E",x"3A",x"0B",x"81",x"0E",x"B0",x"0E",x"3A", -- 0x01F0
    x"0B",x"DD",x"0E",x"13",x"0F",x"3A",x"0B",x"47", -- 0x01F8
    x"0F",x"78",x"0F",x"3A",x"0B",x"A7",x"0F",x"E2", -- 0x0200
    x"0F",x"3A",x"0B",x"74",x"11",x"C7",x"11",x"3A", -- 0x0208
    x"0B",x"F1",x"11",x"17",x"12",x"3A",x"0B",x"18", -- 0x0210
    x"12",x"40",x"12",x"3A",x"0B",x"66",x"12",x"92", -- 0x0218
    x"12",x"3A",x"0B",x"BE",x"12",x"DD",x"12",x"3A", -- 0x0220
    x"0B",x"F6",x"12",x"19",x"13",x"3A",x"0B",x"3A", -- 0x0228
    x"13",x"7A",x"13",x"3A",x"0B",x"B8",x"13",x"EC", -- 0x0230
    x"13",x"3A",x"0B",x"1E",x"14",x"48",x"14",x"3A", -- 0x0238
    x"0B",x"34",x"10",x"CA",x"10",x"3A",x"0B",x"1F", -- 0x0240
    x"0B",x"3F",x"0A",x"5F",x"07",x"91",x"8D",x"8D", -- 0x0248
    x"8D",x"91",x"8D",x"8D",x"8D",x"92",x"92",x"91", -- 0x0250
    x"91",x"AF",x"A0",x"92",x"92",x"91",x"91",x"8F", -- 0x0258
    x"8F",x"96",x"96",x"94",x"92",x"91",x"8F",x"AD", -- 0x0260
    x"A0",x"FF",x"1F",x"05",x"5F",x"07",x"8D",x"91", -- 0x0268
    x"88",x"91",x"8D",x"91",x"88",x"91",x"8F",x"92", -- 0x0270
    x"88",x"92",x"8F",x"92",x"88",x"92",x"8F",x"92", -- 0x0278
    x"88",x"92",x"8F",x"92",x"88",x"92",x"8F",x"92", -- 0x0280
    x"88",x"92",x"B1",x"A0",x"FF",x"1F",x"05",x"5F", -- 0x0288
    x"07",x"80",x"8D",x"80",x"8D",x"80",x"8D",x"80", -- 0x0290
    x"8D",x"80",x"8F",x"80",x"8F",x"80",x"8F",x"80", -- 0x0298
    x"8F",x"80",x"8F",x"80",x"8F",x"80",x"8F",x"80", -- 0x02A0
    x"8F",x"80",x"8F",x"80",x"8F",x"AD",x"A0",x"FF", -- 0x02A8
    x"E7",x"3E",x"01",x"32",x"A3",x"42",x"32",x"A6", -- 0x02B0
    x"42",x"F7",x"C3",x"61",x"09",x"DD",x"21",x"80", -- 0x02B8
    x"42",x"C3",x"A1",x"07",x"E7",x"F7",x"C9",x"DD", -- 0x02C0
    x"21",x"88",x"42",x"C3",x"A1",x"07",x"1F",x"0C", -- 0x02C8
    x"3F",x"0F",x"5F",x"07",x"AD",x"80",x"8A",x"B2", -- 0x02D0
    x"B2",x"B6",x"74",x"72",x"71",x"6F",x"CD",x"AB", -- 0x02D8
    x"AD",x"A8",x"AD",x"AA",x"AD",x"C6",x"FF",x"1F", -- 0x02E0
    x"06",x"5F",x"07",x"AA",x"AD",x"AA",x"AD",x"A6", -- 0x02E8
    x"AD",x"AA",x"AD",x"A8",x"AD",x"AB",x"AD",x"A6", -- 0x02F0
    x"AD",x"CA",x"FF",x"1F",x"0B",x"3F",x"0C",x"5F", -- 0x02F8
    x"07",x"8D",x"8F",x"91",x"92",x"B4",x"B1",x"8D", -- 0x0300
    x"8F",x"91",x"8F",x"AD",x"AD",x"8D",x"8F",x"91", -- 0x0308
    x"92",x"B4",x"B1",x"94",x"92",x"91",x"8F",x"CD", -- 0x0310
    x"FF",x"1F",x"0B",x"5F",x"07",x"85",x"88",x"85", -- 0x0318
    x"88",x"85",x"88",x"85",x"88",x"85",x"88",x"85", -- 0x0320
    x"88",x"85",x"88",x"85",x"88",x"85",x"88",x"85", -- 0x0328
    x"88",x"85",x"88",x"85",x"88",x"86",x"88",x"86", -- 0x0330
    x"88",x"C5",x"FF",x"E7",x"AF",x"32",x"C8",x"42", -- 0x0338
    x"3E",x"02",x"32",x"A3",x"42",x"32",x"A6",x"42", -- 0x0340
    x"F7",x"C3",x"61",x"09",x"DD",x"21",x"80",x"42", -- 0x0348
    x"C3",x"A1",x"07",x"E7",x"F7",x"C9",x"DD",x"21", -- 0x0350
    x"88",x"42",x"C3",x"A1",x"07",x"E7",x"F7",x"C9", -- 0x0358
    x"DD",x"21",x"90",x"42",x"C3",x"A1",x"07",x"E7", -- 0x0360
    x"21",x"A7",x"42",x"34",x"7E",x"FE",x"01",x"28", -- 0x0368
    x"10",x"FE",x"18",x"28",x"11",x"32",x"A3",x"42", -- 0x0370
    x"F7",x"3E",x"01",x"32",x"A5",x"42",x"C3",x"61", -- 0x0378
    x"09",x"36",x"05",x"7E",x"18",x"EF",x"36",x"04", -- 0x0380
    x"3E",x"18",x"18",x"E9",x"E7",x"F7",x"C9",x"DD", -- 0x0388
    x"21",x"80",x"42",x"C3",x"A1",x"07",x"DD",x"21", -- 0x0390
    x"88",x"42",x"C3",x"A1",x"07",x"E7",x"3E",x"03", -- 0x0398
    x"32",x"A3",x"42",x"F7",x"C3",x"5B",x"09",x"3A", -- 0x03A0
    x"A5",x"42",x"A7",x"C2",x"B4",x"07",x"DD",x"21", -- 0x03A8
    x"80",x"42",x"C3",x"A1",x"07",x"1F",x"0B",x"3F", -- 0x03B0
    x"0D",x"5F",x"06",x"9B",x"60",x"7D",x"BB",x"A6", -- 0x03B8
    x"9B",x"60",x"7D",x"BB",x"B8",x"9B",x"60",x"7B", -- 0x03C0
    x"BD",x"80",x"9B",x"99",x"93",x"B8",x"A0",x"8F", -- 0x03C8
    x"60",x"6F",x"8F",x"93",x"B6",x"8F",x"60",x"6F", -- 0x03D0
    x"8F",x"94",x"B8",x"9B",x"60",x"7B",x"BD",x"80", -- 0x03D8
    x"9B",x"99",x"93",x"B4",x"A0",x"FF",x"1F",x"0B", -- 0x03E0
    x"5F",x"06",x"98",x"60",x"77",x"B8",x"B4",x"98", -- 0x03E8
    x"60",x"77",x"B8",x"B4",x"98",x"60",x"76",x"B5", -- 0x03F0
    x"80",x"95",x"96",x"97",x"B4",x"A0",x"8F",x"60", -- 0x03F8
    x"6F",x"8F",x"93",x"B6",x"8F",x"60",x"6D",x"8C", -- 0x0400
    x"8F",x"B4",x"98",x"60",x"76",x"B4",x"80",x"93", -- 0x0408
    x"8F",x"8D",x"AC",x"A0",x"FF",x"1F",x"0B",x"3F", -- 0x0410
    x"0E",x"5F",x"06",x"8F",x"60",x"6F",x"93",x"96", -- 0x0418
    x"BB",x"A0",x"98",x"60",x"78",x"9B",x"98",x"B6", -- 0x0420
    x"A0",x"FF",x"1F",x"0B",x"3F",x"0D",x"5F",x"06", -- 0x0428
    x"8D",x"96",x"B6",x"80",x"97",x"B6",x"94",x"8D", -- 0x0430
    x"B4",x"8D",x"97",x"B7",x"80",x"99",x"B7",x"96", -- 0x0438
    x"8D",x"B6",x"96",x"99",x"B9",x"80",x"9B",x"B9", -- 0x0440
    x"97",x"96",x"94",x"92",x"91",x"94",x"9B",x"99", -- 0x0448
    x"97",x"91",x"D2",x"A0",x"FF",x"1F",x"0B",x"5F", -- 0x0450
    x"06",x"8D",x"92",x"B2",x"80",x"91",x"B2",x"91", -- 0x0458
    x"8D",x"B1",x"8D",x"94",x"B4",x"80",x"96",x"B4", -- 0x0460
    x"92",x"8D",x"B2",x"92",x"96",x"B6",x"80",x"97", -- 0x0468
    x"B6",x"94",x"92",x"91",x"8F",x"8D",x"91",x"97", -- 0x0470
    x"96",x"94",x"8D",x"D2",x"A0",x"FF",x"1F",x"0B", -- 0x0478
    x"3F",x"0D",x"5F",x"06",x"C0",x"A0",x"94",x"60", -- 0x0480
    x"75",x"96",x"9E",x"96",x"9E",x"B6",x"96",x"60", -- 0x0488
    x"75",x"94",x"9D",x"94",x"9D",x"B4",x"9D",x"60", -- 0x0490
    x"73",x"B2",x"BB",x"B9",x"B8",x"B9",x"BB",x"BD", -- 0x0498
    x"94",x"60",x"75",x"96",x"92",x"96",x"92",x"B6", -- 0x04A0
    x"96",x"60",x"79",x"94",x"99",x"94",x"99",x"BD", -- 0x04A8
    x"94",x"60",x"74",x"B4",x"BB",x"B9",x"B8",x"D9", -- 0x04B0
    x"C0",x"FF",x"1F",x"05",x"5F",x"06",x"E0",x"B2", -- 0x04B8
    x"80",x"8D",x"92",x"AD",x"92",x"AD",x"80",x"88", -- 0x04C0
    x"8D",x"A8",x"8D",x"A8",x"80",x"88",x"88",x"A8", -- 0x04C8
    x"88",x"AD",x"80",x"88",x"8D",x"94",x"91",x"8D", -- 0x04D0
    x"B2",x"80",x"8D",x"92",x"AD",x"92",x"AD",x"80", -- 0x04D8
    x"88",x"8D",x"A8",x"8D",x"88",x"94",x"83",x"94", -- 0x04E0
    x"88",x"94",x"88",x"94",x"E0",x"FF",x"1F",x"0B", -- 0x04E8
    x"3F",x"0D",x"5F",x"06",x"B8",x"80",x"96",x"96", -- 0x04F0
    x"94",x"B3",x"B1",x"80",x"AF",x"8D",x"AC",x"CA", -- 0x04F8
    x"AF",x"B6",x"DB",x"9B",x"80",x"8C",x"8D",x"AF", -- 0x0500
    x"B8",x"94",x"80",x"8C",x"8D",x"AF",x"B8",x"94", -- 0x0508
    x"80",x"98",x"99",x"B8",x"B6",x"B8",x"B6",x"D4", -- 0x0510
    x"A0",x"FF",x"1F",x"05",x"5F",x"06",x"A3",x"80", -- 0x0518
    x"AF",x"8F",x"AF",x"A3",x"80",x"AF",x"8F",x"AF", -- 0x0520
    x"A3",x"AF",x"AF",x"AF",x"A3",x"AF",x"8F",x"8F", -- 0x0528
    x"83",x"83",x"A8",x"B4",x"A8",x"B4",x"A8",x"B4", -- 0x0530
    x"A8",x"B4",x"AA",x"B3",x"AF",x"B3",x"B4",x"AF", -- 0x0538
    x"88",x"80",x"FF",x"1F",x"0B",x"3F",x"0D",x"5F", -- 0x0540
    x"06",x"98",x"98",x"98",x"98",x"98",x"98",x"96", -- 0x0548
    x"98",x"99",x"B1",x"80",x"B1",x"B1",x"96",x"96", -- 0x0550
    x"96",x"96",x"B6",x"94",x"96",x"98",x"AF",x"80", -- 0x0558
    x"AF",x"AF",x"98",x"98",x"98",x"98",x"98",x"98", -- 0x0560
    x"96",x"98",x"99",x"99",x"99",x"99",x"B1",x"91", -- 0x0568
    x"94",x"93",x"B3",x"80",x"8F",x"8F",x"98",x"96", -- 0x0570
    x"D4",x"A0",x"FF",x"1F",x"05",x"5F",x"06",x"A8", -- 0x0578
    x"80",x"88",x"C8",x"AA",x"80",x"8A",x"CA",x"AF", -- 0x0580
    x"80",x"8F",x"CF",x"B4",x"80",x"8F",x"AF",x"AC", -- 0x0588
    x"A8",x"80",x"88",x"C8",x"AA",x"80",x"8A",x"CA", -- 0x0590
    x"A3",x"80",x"83",x"C3",x"A8",x"C0",x"FF",x"1F", -- 0x0598
    x"0B",x"3F",x"0D",x"5F",x"06",x"94",x"60",x"72", -- 0x05A0
    x"91",x"94",x"B9",x"9B",x"99",x"96",x"99",x"AF", -- 0x05A8
    x"9B",x"60",x"79",x"98",x"60",x"76",x"94",x"94", -- 0x05B0
    x"96",x"94",x"D4",x"94",x"60",x"72",x"91",x"94", -- 0x05B8
    x"B9",x"9B",x"99",x"96",x"99",x"AF",x"9B",x"60", -- 0x05C0
    x"79",x"98",x"60",x"76",x"94",x"94",x"96",x"98", -- 0x05C8
    x"D9",x"FF",x"1F",x"0B",x"5F",x"06",x"94",x"60", -- 0x05D0
    x"72",x"91",x"94",x"B9",x"98",x"94",x"92",x"91", -- 0x05D8
    x"B2",x"92",x"60",x"76",x"94",x"60",x"74",x"92", -- 0x05E0
    x"92",x"92",x"92",x"D1",x"94",x"60",x"72",x"91", -- 0x05E8
    x"94",x"B9",x"98",x"94",x"92",x"91",x"B2",x"92", -- 0x05F0
    x"60",x"76",x"94",x"60",x"74",x"92",x"92",x"92", -- 0x05F8
    x"92",x"D1",x"FF",x"1F",x"0B",x"3F",x"0D",x"5F", -- 0x0600
    x"06",x"88",x"86",x"65",x"68",x"6D",x"71",x"B4", -- 0x0608
    x"80",x"92",x"71",x"74",x"6D",x"71",x"A8",x"80", -- 0x0610
    x"91",x"6F",x"72",x"6C",x"6F",x"A8",x"80",x"92", -- 0x0618
    x"71",x"74",x"6D",x"71",x"A8",x"88",x"60",x"66", -- 0x0620
    x"65",x"68",x"6D",x"71",x"B4",x"8D",x"60",x"6B", -- 0x0628
    x"6A",x"6D",x"72",x"76",x"B9",x"98",x"96",x"94", -- 0x0630
    x"60",x"71",x"96",x"60",x"71",x"94",x"60",x"71", -- 0x0638
    x"72",x"68",x"6C",x"6F",x"B4",x"80",x"92",x"71", -- 0x0640
    x"68",x"6D",x"71",x"B4",x"80",x"91",x"6F",x"68", -- 0x0648
    x"71",x"60",x"6F",x"68",x"71",x"60",x"6F",x"68", -- 0x0650
    x"74",x"60",x"D9",x"FF",x"1F",x"0B",x"5F",x"06", -- 0x0658
    x"A0",x"AD",x"AC",x"A0",x"AA",x"A8",x"A0",x"A6", -- 0x0660
    x"A5",x"A0",x"A8",x"A6",x"A0",x"AD",x"A7",x"A0", -- 0x0668
    x"AA",x"A8",x"A0",x"A5",x"A6",x"A5",x"A8",x"A6", -- 0x0670
    x"A0",x"A8",x"A5",x"A0",x"A6",x"A8",x"A6",x"C5", -- 0x0678
    x"FF",x"1F",x"0B",x"3F",x"0D",x"5F",x"06",x"94", -- 0x0680
    x"99",x"99",x"9B",x"9B",x"9D",x"9D",x"98",x"9B", -- 0x0688
    x"B9",x"B6",x"B4",x"80",x"92",x"91",x"8F",x"91", -- 0x0690
    x"92",x"94",x"B4",x"99",x"98",x"94",x"96",x"98", -- 0x0698
    x"B9",x"80",x"92",x"91",x"8F",x"91",x"92",x"94", -- 0x06A0
    x"B4",x"99",x"98",x"94",x"96",x"98",x"B9",x"FF", -- 0x06A8
    x"1F",x"0B",x"5F",x"06",x"94",x"94",x"94",x"94", -- 0x06B0
    x"94",x"94",x"94",x"92",x"92",x"B1",x"B3",x"B4", -- 0x06B8
    x"80",x"8F",x"8D",x"8C",x"8D",x"8F",x"8F",x"8F", -- 0x06C0
    x"B4",x"92",x"92",x"92",x"92",x"B1",x"80",x"8F", -- 0x06C8
    x"8D",x"8C",x"8D",x"8F",x"8F",x"8F",x"B4",x"92", -- 0x06D0
    x"92",x"92",x"92",x"B1",x"FF",x"1F",x"0B",x"3F", -- 0x06D8
    x"0D",x"5F",x"06",x"87",x"60",x"68",x"AA",x"80", -- 0x06E0
    x"8F",x"8E",x"60",x"6C",x"CA",x"8F",x"60",x"6F", -- 0x06E8
    x"6E",x"71",x"94",x"9A",x"60",x"78",x"96",x"8E", -- 0x06F0
    x"8F",x"93",x"8A",x"80",x"87",x"60",x"68",x"AA", -- 0x06F8
    x"80",x"8F",x"8E",x"60",x"6C",x"CA",x"8F",x"60", -- 0x0700
    x"6F",x"6E",x"71",x"94",x"9A",x"60",x"78",x"96", -- 0x0708
    x"8E",x"CF",x"FF",x"1F",x"0B",x"5F",x"06",x"87", -- 0x0710
    x"60",x"68",x"AA",x"80",x"8F",x"8E",x"60",x"6C", -- 0x0718
    x"CA",x"8F",x"60",x"6F",x"6E",x"6E",x"91",x"96", -- 0x0720
    x"60",x"74",x"91",x"88",x"87",x"88",x"87",x"80", -- 0x0728
    x"87",x"60",x"68",x"AA",x"80",x"87",x"88",x"60", -- 0x0730
    x"68",x"C7",x"8F",x"60",x"6F",x"6E",x"6E",x"91", -- 0x0738
    x"96",x"60",x"74",x"91",x"88",x"C7",x"FF",x"1F", -- 0x0740
    x"0B",x"3F",x"0D",x"5F",x"06",x"8A",x"8F",x"8E", -- 0x0748
    x"91",x"AA",x"8C",x"8E",x"8F",x"93",x"AA",x"8A", -- 0x0750
    x"8F",x"8E",x"91",x"AA",x"8C",x"8E",x"8F",x"93", -- 0x0758
    x"AA",x"87",x"60",x"68",x"AA",x"80",x"8F",x"8E", -- 0x0760
    x"60",x"6C",x"CA",x"8F",x"60",x"6F",x"6E",x"71", -- 0x0768
    x"94",x"9A",x"60",x"78",x"96",x"8E",x"CF",x"FF", -- 0x0770
    x"1F",x"0B",x"5F",x"06",x"8A",x"87",x"88",x"88", -- 0x0778
    x"A8",x"88",x"88",x"87",x"8A",x"A7",x"87",x"87", -- 0x0780
    x"88",x"88",x"A8",x"88",x"88",x"87",x"8A",x"A7", -- 0x0788
    x"87",x"60",x"68",x"AA",x"80",x"87",x"88",x"60", -- 0x0790
    x"68",x"C7",x"8F",x"60",x"6F",x"6E",x"6E",x"91", -- 0x0798
    x"96",x"60",x"74",x"91",x"88",x"C7",x"FF",x"1F", -- 0x07A0
    x"0B",x"3F",x"0C",x"5F",x"06",x"B4",x"91",x"8D", -- 0x07A8
    x"B9",x"98",x"96",x"B4",x"99",x"91",x"8F",x"B4", -- 0x07B0
    x"80",x"94",x"94",x"94",x"94",x"96",x"94",x"91", -- 0x07B8
    x"8D",x"99",x"99",x"99",x"99",x"9B",x"99",x"96", -- 0x07C0
    x"92",x"94",x"94",x"94",x"94",x"96",x"94",x"91", -- 0x07C8
    x"8D",x"99",x"99",x"99",x"99",x"9B",x"99",x"96", -- 0x07D0
    x"92",x"94",x"91",x"80",x"91",x"B9",x"B1",x"94", -- 0x07D8
    x"CF",x"FF",x"1F",x"05",x"5F",x"06",x"D9",x"D6", -- 0x07E0
    x"D9",x"D8",x"8D",x"91",x"88",x"91",x"8D",x"91", -- 0x07E8
    x"88",x"91",x"8D",x"92",x"8A",x"92",x"8D",x"92", -- 0x07F0
    x"8A",x"92",x"8D",x"91",x"88",x"91",x"8D",x"91"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
