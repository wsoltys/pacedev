-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_SND_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_SND_0 is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"05",x"00",x"22",x"00",x"40",x"C3",x"0B",x"02", -- 0x0000
    x"D3",x"80",x"78",x"D3",x"40",x"CA",x"FF",x"FF", -- 0x0008
    x"C3",x"B7",x"01",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0010
    x"C3",x"7C",x"01",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0018
    x"C3",x"C7",x"01",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0020
    x"C3",x"3C",x"01",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0028
    x"C3",x"60",x"01",x"3D",x"FF",x"CA",x"FF",x"FF", -- 0x0030
    x"08",x"DA",x"22",x"6E",x"00",x"E6",x"3D",x"0D", -- 0x0038
    x"CE",x"C2",x"01",x"B7",x"28",x"2B",x"57",x"FD", -- 0x0040
    x"FF",x"20",x"02",x"C7",x"E5",x"0F",x"4F",x"79", -- 0x0048
    x"AA",x"28",x"07",x"7A",x"B7",x"28",x"03",x"79", -- 0x0050
    x"18",x"3E",x"79",x"E5",x"0F",x"20",x"38",x"79", -- 0x0058
    x"C5",x"11",x"07",x"07",x"07",x"CB",x"7F",x"28", -- 0x0060
    x"2D",x"CB",x"BF",x"18",x"13",x"DA",x"08",x"FB", -- 0x0068
    x"CA",x"05",x"05",x"22",x"40",x"40",x"77",x"23", -- 0x0070
    x"10",x"FC",x"3D",x"07",x"05",x"3F",x"CF",x"CA", -- 0x0078
    x"CE",x"E5",x"00",x"D0",x"CE",x"8C",x"00",x"AF", -- 0x0080
    x"77",x"23",x"77",x"CA",x"47",x"22",x"3D",x"40", -- 0x0088
    x"12",x"01",x"00",x"1A",x"10",x"FE",x"CA",x"31", -- 0x0090
    x"45",x"40",x"CE",x"E5",x"00",x"D8",x"CE",x"E5", -- 0x0098
    x"00",x"38",x"38",x"39",x"40",x"40",x"CE",x"01", -- 0x00A0
    x"02",x"47",x"39",x"41",x"40",x"CE",x"01",x"02", -- 0x00A8
    x"4F",x"39",x"44",x"40",x"CE",x"01",x"02",x"31", -- 0x00B0
    x"4A",x"40",x"39",x"45",x"40",x"CE",x"01",x"02", -- 0x00B8
    x"5F",x"22",x"4A",x"40",x"55",x"78",x"BA",x"38", -- 0x00C0
    x"02",x"7A",x"B9",x"38",x"02",x"79",x"BB",x"D0", -- 0x00C8
    x"1D",x"02",x"B8",x"28",x"06",x"1C",x"BA",x"28", -- 0x00D0
    x"02",x"1C",x"7B",x"CE",x"8C",x"00",x"39",x"45", -- 0x00D8
    x"40",x"77",x"23",x"35",x"00",x"CA",x"0D",x"02", -- 0x00E0
    x"22",x"40",x"40",x"BD",x"28",x"0D",x"0C",x"23", -- 0x00E8
    x"23",x"BD",x"28",x"08",x"0C",x"23",x"23",x"BD", -- 0x00F0
    x"28",x"01",x"AF",x"CA",x"23",x"35",x"00",x"7A", -- 0x00F8
    x"37",x"CA",x"22",x"83",x"01",x"5F",x"15",x"00", -- 0x0100
    x"1A",x"7D",x"CA",x"70",x"23",x"7C",x"D5",x"44", -- 0x0108
    x"20",x"FA",x"FA",x"3E",x"31",x"80",x"41",x"EE", -- 0x0110
    x"55",x"12",x"3F",x"00",x"CE",x"6E",x"01",x"3D", -- 0x0118
    x"08",x"05",x"00",x"CF",x"3D",x"0A",x"CF",x"3D", -- 0x0120
    x"09",x"CF",x"3D",x"07",x"05",x"3F",x"CF",x"22", -- 0x0128
    x"00",x"60",x"21",x"4D",x"40",x"77",x"FB",x"22", -- 0x0130
    x"3F",x"40",x"34",x"3D",x"0F",x"CE",x"C2",x"01", -- 0x0138
    x"E5",x"08",x"20",x"F7",x"3D",x"0F",x"CE",x"C2", -- 0x0140
    x"01",x"E5",x"08",x"28",x"F7",x"F3",x"3D",x"02", -- 0x0148
    x"31",x"4B",x"40",x"22",x"42",x"40",x"7D",x"2B", -- 0x0150
    x"B7",x"28",x"30",x"7D",x"CE",x"E8",x"02",x"FB", -- 0x0158
    x"00",x"00",x"00",x"F3",x"22",x"4B",x"40",x"34", -- 0x0160
    x"22",x"43",x"40",x"7D",x"2B",x"B7",x"28",x"22", -- 0x0168
    x"7D",x"CE",x"E8",x"02",x"FB",x"00",x"00",x"00", -- 0x0170
    x"F3",x"22",x"4B",x"40",x"34",x"22",x"46",x"40", -- 0x0178
    x"7D",x"2B",x"B7",x"28",x"11",x"7D",x"CE",x"E8", -- 0x0180
    x"02",x"18",x"AB",x"7D",x"CE",x"DA",x"02",x"18", -- 0x0188
    x"CD",x"7D",x"CE",x"DA",x"02",x"18",x"DE",x"7D", -- 0x0190
    x"CE",x"DA",x"02",x"18",x"9A",x"87",x"5F",x"15", -- 0x0198
    x"00",x"1A",x"5D",x"23",x"55",x"EB",x"EA",x"9C", -- 0x01A0
    x"01",x"0F",x"03",x"BE",x"03",x"5E",x"04",x"81", -- 0x01A8
    x"14",x"66",x"14",x"9E",x"0B",x"8E",x"04",x"67", -- 0x01B0
    x"0B",x"7F",x"07",x"8B",x"07",x"8D",x"07",x"B0", -- 0x01B8
    x"09",x"C4",x"09",x"8C",x"0B",x"16",x"10",x"EB", -- 0x01C0
    x"05",x"3B",x"0B",x"53",x"0B",x"5E",x"0B",x"00", -- 0x01C8
    x"00",x"06",x"06",x"23",x"10",x"C3",x"06",x"3E", -- 0x01D0
    x"05",x"22",x"A7",x"02",x"CE",x"9E",x"02",x"39", -- 0x01D8
    x"4B",x"40",x"CE",x"8C",x"00",x"23",x"77",x"CA", -- 0x01E0
    x"B7",x"C8",x"22",x"26",x"01",x"E6",x"22",x"F3", -- 0x01E8
    x"02",x"18",x"A9",x"33",x"00",x"33",x"03",x"D1", -- 0x01F0
    x"03",x"76",x"04",x"8C",x"14",x"71",x"14",x"A7", -- 0x01F8
    x"0B",x"A9",x"04",x"8F",x"0B",x"92",x"07",x"97", -- 0x0200
    x"07",x"9E",x"07",x"BE",x"09",x"C7",x"09",x"95", -- 0x0208
    x"0B",x"25",x"10",x"0D",x"07",x"4C",x"0B",x"55", -- 0x0210
    x"0B",x"60",x"0B",x"00",x"00",x"1C",x"06",x"2E", -- 0x0218
    x"10",x"E6",x"06",x"62",x"05",x"B7",x"C8",x"CE", -- 0x0220
    x"9C",x"01",x"39",x"4B",x"40",x"C3",x"84",x"00", -- 0x0228
    x"39",x"4B",x"40",x"E5",x"03",x"C8",x"C5",x"07", -- 0x0230
    x"05",x"00",x"CF",x"CA",x"39",x"4B",x"40",x"3E", -- 0x0238
    x"87",x"47",x"CE",x"0A",x"03",x"04",x"78",x"D3", -- 0x0240
    x"80",x"7C",x"D3",x"40",x"CA",x"39",x"4B",x"40", -- 0x0248
    x"3E",x"87",x"47",x"D3",x"80",x"DB",x"40",x"6F", -- 0x0250
    x"04",x"78",x"D3",x"80",x"DB",x"40",x"67",x"CA", -- 0x0258
    x"12",x"04",x"7F",x"39",x"4B",x"40",x"47",x"CB", -- 0x0260
    x"01",x"CB",x"03",x"10",x"F9",x"3D",x"07",x"D3", -- 0x0268
    x"80",x"39",x"4C",x"40",x"A1",x"B3",x"31",x"4C", -- 0x0270
    x"40",x"D3",x"40",x"CA",x"39",x"4B",x"40",x"C5", -- 0x0278
    x"07",x"CF",x"CA",x"00",x"06",x"09",x"0E",x"18", -- 0x0280
    x"07",x"0D",x"0C",x"05",x"16",x"14",x"13",x"10", -- 0x0288
    x"0F",x"04",x"15",x"03",x"11",x"12",x"01",x"0A", -- 0x0290
    x"08",x"02",x"15",x"17",x"39",x"4B",x"40",x"47", -- 0x0298
    x"3D",x"84",x"07",x"10",x"FE",x"5F",x"15",x"FF", -- 0x02A0
    x"CE",x"6E",x"01",x"CE",x"30",x"01",x"18",x"17", -- 0x02A8
    x"12",x"80",x"FB",x"18",x"AD",x"CF",x"CA",x"39", -- 0x02B0
    x"4B",x"40",x"E5",x"03",x"C8",x"C5",x"07",x"18", -- 0x02B8
    x"00",x"D3",x"80",x"DB",x"40",x"47",x"CA",x"02", -- 0x02C0
    x"00",x"00",x"12",x"FF",x"FC",x"39",x"4B",x"40", -- 0x02C8
    x"FD",x"01",x"28",x"16",x"38",x"08",x"15",x"F3", -- 0x02D0
    x"CB",x"00",x"CB",x"00",x"18",x"0B",x"12",x"3F", -- 0x02D8
    x"FF",x"CB",x"38",x"CB",x"1A",x"CB",x"38",x"CB", -- 0x02E0
    x"1A",x"29",x"4D",x"40",x"7C",x"A1",x"B0",x"67", -- 0x02E8
    x"7E",x"A3",x"B2",x"6F",x"21",x"4D",x"40",x"77", -- 0x02F0
    x"CA",x"02",x"00",x"03",x"C3",x"C9",x"01",x"02", -- 0x02F8
    x"00",x"02",x"18",x"C5",x"02",x"00",x"01",x"18", -- 0x0300
    x"C2",x"D3",x"80",x"7E",x"D3",x"40",x"CA",x"E7", -- 0x0308
    x"3D",x"20",x"22",x"60",x"40",x"77",x"3D",x"03", -- 0x0310
    x"23",x"77",x"3D",x"14",x"23",x"77",x"3D",x"02", -- 0x0318
    x"23",x"77",x"AF",x"23",x"77",x"22",x"10",x"00", -- 0x0320
    x"21",x"66",x"40",x"2D",x"20",x"EF",x"F7",x"05", -- 0x0328
    x"0A",x"DF",x"CA",x"39",x"64",x"40",x"A7",x"28", -- 0x0330
    x"0E",x"FD",x"02",x"28",x"1F",x"FD",x"03",x"38", -- 0x0338
    x"2B",x"28",x"4A",x"C3",x"72",x"05",x"22",x"60", -- 0x0340
    x"40",x"36",x"20",x"6F",x"35",x"20",x"D7",x"3E", -- 0x0348
    x"28",x"04",x"47",x"DF",x"18",x"66",x"22",x"64", -- 0x0350
    x"40",x"34",x"18",x"F5",x"22",x"00",x"03",x"21", -- 0x0358
    x"67",x"40",x"EF",x"05",x"08",x"DF",x"22",x"64", -- 0x0360
    x"40",x"34",x"18",x"4F",x"22",x"62",x"40",x"36", -- 0x0368
    x"20",x"4A",x"35",x"03",x"CE",x"4E",x"01",x"B7", -- 0x0370
    x"12",x"08",x"00",x"EE",x"51",x"EF",x"22",x"61", -- 0x0378
    x"40",x"36",x"20",x"37",x"35",x"14",x"22",x"64", -- 0x0380
    x"40",x"34",x"18",x"2F",x"22",x"63",x"40",x"36", -- 0x0388
    x"20",x"1E",x"35",x"02",x"B7",x"29",x"67",x"40", -- 0x0390
    x"12",x"20",x"00",x"EE",x"51",x"21",x"67",x"40", -- 0x0398
    x"EF",x"29",x"66",x"40",x"2B",x"7E",x"B4",x"20", -- 0x03A0
    x"0B",x"22",x"64",x"40",x"34",x"18",x"0C",x"29", -- 0x03A8
    x"67",x"40",x"18",x"EC",x"21",x"66",x"40",x"22", -- 0x03B0
    x"64",x"40",x"36",x"AF",x"CA",x"3D",x"80",x"31", -- 0x03B8
    x"5E",x"40",x"05",x"0D",x"CE",x"7C",x"01",x"22", -- 0x03C0
    x"70",x"00",x"CE",x"3C",x"01",x"F7",x"CE",x"04", -- 0x03C8
    x"03",x"CA",x"39",x"5E",x"40",x"3E",x"31",x"5E", -- 0x03D0
    x"40",x"28",x"26",x"FD",x"FF",x"28",x"39",x"FD", -- 0x03D8
    x"20",x"38",x"09",x"FD",x"30",x"38",x"0C",x"FD", -- 0x03E0
    x"70",x"38",x"01",x"AF",x"CA",x"05",x"00",x"CE", -- 0x03E8
    x"7C",x"01",x"CA",x"22",x"3C",x"00",x"CE",x"3C", -- 0x03F0
    x"01",x"05",x"0B",x"CE",x"7C",x"01",x"AF",x"CA", -- 0x03F8
    x"CE",x"04",x"03",x"3D",x"80",x"31",x"5D",x"40", -- 0x0400
    x"05",x"09",x"CE",x"7C",x"01",x"22",x"FC",x"00", -- 0x0408
    x"CE",x"3C",x"01",x"F7",x"AF",x"31",x"5E",x"40", -- 0x0410
    x"CA",x"39",x"5D",x"40",x"3E",x"31",x"5D",x"40", -- 0x0418
    x"FD",x"42",x"38",x"0B",x"CE",x"4E",x"01",x"2E", -- 0x0420
    x"2E",x"EF",x"AF",x"31",x"5E",x"40",x"CA",x"FD", -- 0x0428
    x"40",x"28",x"0D",x"B7",x"28",x"12",x"CE",x"4E", -- 0x0430
    x"01",x"2C",x"2C",x"EF",x"AF",x"31",x"5E",x"40", -- 0x0438
    x"CA",x"D7",x"06",x"DF",x"C3",x"33",x"04",x"D7", -- 0x0440
    x"06",x"28",x"0F",x"DF",x"22",x"00",x"00",x"CE", -- 0x0448
    x"3C",x"01",x"3D",x"80",x"31",x"5D",x"40",x"C3", -- 0x0450
    x"1A",x"04",x"3D",x"FF",x"CA",x"CE",x"C7",x"01", -- 0x0458
    x"CE",x"60",x"01",x"22",x"00",x"02",x"CE",x"3C", -- 0x0460
    x"01",x"05",x"09",x"CE",x"7C",x"01",x"22",x"90", -- 0x0468
    x"01",x"21",x"30",x"42",x"CA",x"29",x"30",x"42", -- 0x0470
    x"2B",x"21",x"30",x"42",x"7C",x"B6",x"3D",x"FF", -- 0x0478
    x"C8",x"CE",x"4E",x"01",x"12",x"03",x"00",x"1A", -- 0x0480
    x"CE",x"3C",x"01",x"AF",x"CA",x"E7",x"3D",x"08", -- 0x0488
    x"31",x"70",x"42",x"3D",x"0C",x"31",x"72",x"42", -- 0x0490
    x"3D",x"10",x"31",x"71",x"42",x"AF",x"31",x"73", -- 0x0498
    x"42",x"22",x"50",x"00",x"EF",x"F7",x"05",x"00", -- 0x04A0
    x"DF",x"CA",x"39",x"73",x"42",x"A7",x"28",x"17", -- 0x04A8
    x"FD",x"02",x"28",x"22",x"FD",x"03",x"38",x"21", -- 0x04B0
    x"28",x"2C",x"22",x"71",x"42",x"36",x"3D",x"FF", -- 0x04B8
    x"C8",x"AF",x"31",x"73",x"42",x"AF",x"CA",x"D7", -- 0x04C0
    x"3C",x"FD",x"0E",x"20",x"04",x"22",x"73",x"42", -- 0x04C8
    x"34",x"47",x"DF",x"18",x"F0",x"CE",x"EB",x"04", -- 0x04D0
    x"18",x"EB",x"D7",x"3E",x"20",x"04",x"22",x"73", -- 0x04D8
    x"42",x"34",x"47",x"DF",x"18",x"DF",x"CE",x"F8", -- 0x04E0
    x"04",x"18",x"D9",x"22",x"70",x"42",x"36",x"C0", -- 0x04E8
    x"3D",x"08",x"77",x"22",x"73",x"42",x"34",x"CA", -- 0x04F0
    x"22",x"72",x"42",x"36",x"C0",x"3D",x"0C",x"77", -- 0x04F8
    x"22",x"73",x"42",x"34",x"CA",x"CE",x"04",x"03", -- 0x0500
    x"22",x"00",x"02",x"21",x"75",x"42",x"F7",x"05", -- 0x0508
    x"05",x"DF",x"3D",x"08",x"31",x"76",x"42",x"AF", -- 0x0510
    x"31",x"78",x"42",x"CA",x"39",x"78",x"42",x"FD", -- 0x0518
    x"02",x"28",x"34",x"FD",x"01",x"28",x"48",x"FD", -- 0x0520
    x"03",x"28",x"6A",x"FD",x"04",x"28",x"75",x"22", -- 0x0528
    x"76",x"42",x"36",x"20",x"15",x"35",x"08",x"12", -- 0x0530
    x"F0",x"FF",x"29",x"75",x"42",x"1A",x"21",x"75", -- 0x0538
    x"42",x"7C",x"A7",x"20",x"06",x"7E",x"FD",x"38", -- 0x0540
    x"38",x"03",x"EF",x"AF",x"CA",x"3D",x"20",x"31", -- 0x0548
    x"76",x"42",x"44",x"3D",x"02",x"18",x"11",x"22", -- 0x0550
    x"76",x"42",x"36",x"20",x"ED",x"35",x"06",x"3D", -- 0x0558
    x"03",x"22",x"60",x"00",x"05",x"01",x"21",x"75", -- 0x0560
    x"42",x"31",x"78",x"42",x"DF",x"AF",x"CA",x"22", -- 0x0568
    x"76",x"42",x"36",x"20",x"D5",x"35",x"05",x"12", -- 0x0570
    x"FC",x"FF",x"29",x"75",x"42",x"1A",x"21",x"75", -- 0x0578
    x"42",x"7C",x"A7",x"20",x"C6",x"7E",x"FD",x"30", -- 0x0580
    x"30",x"C0",x"3D",x"30",x"31",x"76",x"42",x"44", -- 0x0588
    x"3D",x"03",x"18",x"D6",x"22",x"76",x"42",x"36", -- 0x0590
    x"20",x"B2",x"35",x"04",x"3D",x"04",x"22",x"60", -- 0x0598
    x"00",x"05",x"04",x"18",x"C2",x"22",x"76",x"42", -- 0x05A0
    x"36",x"20",x"A0",x"35",x"04",x"12",x"10",x"00", -- 0x05A8
    x"29",x"75",x"42",x"1A",x"21",x"75",x"42",x"7C", -- 0x05B0
    x"A7",x"28",x"8F",x"7E",x"FD",x"80",x"38",x"89", -- 0x05B8
    x"C3",x"06",x"06",x"AF",x"22",x"10",x"42",x"77", -- 0x05C0
    x"23",x"35",x"04",x"23",x"35",x"04",x"23",x"35", -- 0x05C8
    x"04",x"23",x"35",x"68",x"CE",x"B0",x"01",x"3D", -- 0x05D0
    x"05",x"05",x"18",x"CF",x"05",x"04",x"CE",x"7C", -- 0x05D8
    x"01",x"CE",x"C7",x"01",x"CA",x"CE",x"1C",x"05", -- 0x05E0
    x"CE",x"EE",x"06",x"AF",x"CA",x"39",x"10",x"42", -- 0x05E8
    x"CB",x"47",x"28",x"10",x"22",x"11",x"42",x"36", -- 0x05F0
    x"C0",x"35",x"04",x"05",x"00",x"CE",x"7C",x"01", -- 0x05F8
    x"0D",x"02",x"18",x"10",x"22",x"12",x"42",x"36", -- 0x0600
    x"C0",x"35",x"04",x"39",x"13",x"42",x"47",x"CE", -- 0x0608
    x"7C",x"01",x"0D",x"02",x"39",x"10",x"42",x"AA", -- 0x0610
    x"31",x"10",x"42",x"CA",x"22",x"14",x"42",x"36", -- 0x0618
    x"C0",x"35",x"68",x"22",x"13",x"42",x"39",x"10", -- 0x0620
    x"42",x"CB",x"4F",x"20",x"0A",x"34",x"3D",x"07", -- 0x0628
    x"BD",x"0D",x"01",x"28",x"DF",x"CA",x"36",x"7D", -- 0x0630
    x"3C",x"C0",x"E2",x"3E",x"CA",x"E7",x"3D",x"20", -- 0x0638
    x"22",x"E0",x"42",x"77",x"3D",x"03",x"23",x"77", -- 0x0640
    x"3D",x"14",x"23",x"77",x"3D",x"02",x"23",x"77", -- 0x0648
    x"23",x"35",x"00",x"22",x"10",x"00",x"21",x"E6", -- 0x0650
    x"42",x"2D",x"20",x"EF",x"F7",x"05",x"0A",x"DF", -- 0x0658
    x"CA",x"39",x"E4",x"42",x"A7",x"28",x"1C",x"FD", -- 0x0660
    x"02",x"28",x"1F",x"FD",x"03",x"38",x"2B",x"28", -- 0x0668
    x"4A",x"D7",x"3E",x"28",x"04",x"47",x"DF",x"AF", -- 0x0670
    x"CA",x"AF",x"31",x"A6",x"41",x"3E",x"CA",x"47", -- 0x0678
    x"DF",x"18",x"65",x"22",x"E4",x"42",x"34",x"AF", -- 0x0680
    x"18",x"F6",x"22",x"00",x"03",x"21",x"E7",x"42", -- 0x0688
    x"EF",x"05",x"08",x"DF",x"22",x"E4",x"42",x"34", -- 0x0690
    x"18",x"4F",x"22",x"E2",x"42",x"36",x"20",x"4A", -- 0x0698
    x"35",x"03",x"CE",x"4E",x"01",x"B7",x"12",x"08", -- 0x06A0
    x"00",x"EE",x"51",x"EF",x"22",x"E1",x"42",x"36", -- 0x06A8
    x"20",x"37",x"35",x"14",x"22",x"E4",x"42",x"34", -- 0x06B0
    x"18",x"2F",x"22",x"E3",x"42",x"36",x"20",x"1E", -- 0x06B8
    x"35",x"02",x"B7",x"29",x"E7",x"42",x"12",x"20", -- 0x06C0
    x"00",x"EE",x"51",x"21",x"E7",x"42",x"EF",x"29", -- 0x06C8
    x"E6",x"42",x"2B",x"7E",x"B4",x"20",x"0B",x"22", -- 0x06D0
    x"E4",x"42",x"34",x"18",x"0C",x"29",x"E7",x"42", -- 0x06D8
    x"18",x"EC",x"21",x"E6",x"42",x"22",x"E4",x"42", -- 0x06E0
    x"36",x"AF",x"CA",x"22",x"50",x"00",x"21",x"80", -- 0x06E8
    x"42",x"22",x"24",x"0A",x"21",x"81",x"42",x"3D", -- 0x06F0
    x"00",x"31",x"84",x"42",x"05",x"0E",x"CE",x"7C", -- 0x06F8
    x"01",x"22",x"50",x"00",x"CE",x"3C",x"01",x"CE", -- 0x0700
    x"60",x"01",x"CE",x"C7",x"01",x"CA",x"29",x"80", -- 0x0708
    x"42",x"2B",x"21",x"80",x"42",x"7C",x"B6",x"3D", -- 0x0710
    x"00",x"28",x"47",x"39",x"84",x"42",x"CB",x"47", -- 0x0718
    x"3D",x"00",x"28",x"0D",x"22",x"81",x"42",x"36", -- 0x0720
    x"C0",x"35",x"24",x"05",x"0E",x"CE",x"7C",x"01", -- 0x0728
    x"18",x"26",x"CE",x"4E",x"01",x"12",x"09",x"00", -- 0x0730
    x"39",x"84",x"42",x"CB",x"4F",x"28",x"04",x"AF", -- 0x0738
    x"EE",x"51",x"3D",x"1A",x"CE",x"3C",x"01",x"0D", -- 0x0740
    x"01",x"CE",x"5A",x"07",x"22",x"83",x"42",x"36", -- 0x0748
    x"C0",x"35",x"0A",x"47",x"CE",x"7C",x"01",x"0D", -- 0x0750
    x"02",x"39",x"84",x"42",x"AA",x"31",x"84",x"42", -- 0x0758
    x"AF",x"CA",x"22",x"84",x"42",x"CB",x"55",x"20", -- 0x0760
    x"0D",x"CE",x"EB",x"05",x"05",x"00",x"CE",x"7C", -- 0x0768
    x"01",x"22",x"84",x"42",x"CB",x"D5",x"CA",x"05", -- 0x0770
    x"00",x"CE",x"7C",x"01",x"3D",x"FF",x"CA",x"E7", -- 0x0778
    x"AF",x"31",x"C8",x"41",x"31",x"A3",x"41",x"F7", -- 0x0780
    x"C3",x"62",x"0A",x"E7",x"F7",x"CA",x"E7",x"F7", -- 0x0788
    x"CA",x"DE",x"22",x"80",x"41",x"18",x"09",x"DE", -- 0x0790
    x"22",x"88",x"41",x"18",x"04",x"DE",x"22",x"90", -- 0x0798
    x"41",x"DE",x"7D",x"00",x"FD",x"FF",x"28",x"06", -- 0x07A0
    x"CE",x"B7",x"07",x"AF",x"CA",x"AF",x"31",x"A6", -- 0x07A8
    x"41",x"31",x"A5",x"41",x"3D",x"FF",x"CA",x"DE", -- 0x07B0
    x"36",x"02",x"C0",x"39",x"A1",x"41",x"DE",x"77", -- 0x07B8
    x"02",x"DE",x"CB",x"00",x"45",x"C1",x"D6",x"07", -- 0x07C0
    x"DE",x"7D",x"07",x"D5",x"02",x"F9",x"D6",x"07", -- 0x07C8
    x"DE",x"77",x"07",x"47",x"DF",x"DE",x"36",x"00", -- 0x07D0
    x"C0",x"DE",x"6D",x"01",x"DE",x"65",x"03",x"7D", -- 0x07D8
    x"47",x"E5",x"1F",x"C9",x"69",x"08",x"FD",x"1F", -- 0x07E0
    x"C1",x"84",x"08",x"23",x"DE",x"76",x"01",x"DE", -- 0x07E8
    x"74",x"03",x"78",x"E5",x"E0",x"0F",x"0F",x"0F", -- 0x07F0
    x"0F",x"4F",x"05",x"00",x"22",x"06",x"08",x"0A"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
