-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_SND_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_SND_0 is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"C3",x"72",x"02",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0000
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0008
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0010
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0018
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0020
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0028
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0030
    x"08",x"D9",x"3E",x"0E",x"D3",x"40",x"DB",x"80", -- 0x0038
    x"B7",x"28",x"13",x"FE",x"30",x"FA",x"64",x"00", -- 0x0040
    x"FE",x"40",x"F2",x"6B",x"00",x"D6",x"10",x"CD", -- 0x0048
    x"6F",x"00",x"D9",x"08",x"FB",x"C9",x"06",x"0C", -- 0x0050
    x"21",x"00",x"80",x"77",x"23",x"05",x"20",x"FB", -- 0x0058
    x"D9",x"08",x"FB",x"C9",x"CD",x"E7",x"00",x"D9", -- 0x0060
    x"08",x"FB",x"C9",x"D9",x"08",x"FB",x"C9",x"CD", -- 0x0068
    x"A6",x"00",x"B7",x"C8",x"FE",x"01",x"28",x"15", -- 0x0070
    x"FE",x"02",x"28",x"16",x"FE",x"03",x"28",x"17", -- 0x0078
    x"FE",x"04",x"28",x"18",x"FE",x"05",x"28",x"19", -- 0x0080
    x"AF",x"32",x"0A",x"80",x"C9",x"AF",x"32",x"00", -- 0x0088
    x"80",x"C9",x"AF",x"32",x"02",x"80",x"C9",x"AF", -- 0x0090
    x"32",x"04",x"80",x"C9",x"AF",x"32",x"06",x"80", -- 0x0098
    x"C9",x"AF",x"32",x"08",x"80",x"C9",x"06",x"00", -- 0x00A0
    x"21",x"00",x"80",x"BE",x"28",x"1B",x"23",x"23", -- 0x00A8
    x"BE",x"28",x"1B",x"23",x"23",x"BE",x"28",x"1B", -- 0x00B0
    x"23",x"23",x"BE",x"28",x"1B",x"23",x"23",x"BE", -- 0x00B8
    x"28",x"1B",x"23",x"23",x"BE",x"28",x"1B",x"AF", -- 0x00C0
    x"C9",x"23",x"70",x"3E",x"01",x"C9",x"23",x"70", -- 0x00C8
    x"3E",x"02",x"C9",x"23",x"70",x"3E",x"03",x"C9", -- 0x00D0
    x"23",x"70",x"3E",x"04",x"C9",x"23",x"70",x"3E", -- 0x00D8
    x"05",x"C9",x"23",x"70",x"3E",x"06",x"C9",x"32", -- 0x00E0
    x"1A",x"80",x"CD",x"A6",x"00",x"B7",x"C0",x"AF", -- 0x00E8
    x"CD",x"A6",x"00",x"B7",x"20",x"73",x"3A",x"00", -- 0x00F0
    x"80",x"CD",x"F1",x"01",x"32",x"12",x"80",x"3A", -- 0x00F8
    x"02",x"80",x"CD",x"F1",x"01",x"32",x"13",x"80", -- 0x0100
    x"3A",x"04",x"80",x"CD",x"F1",x"01",x"32",x"14", -- 0x0108
    x"80",x"3A",x"1A",x"80",x"CD",x"F1",x"01",x"32", -- 0x0110
    x"15",x"80",x"CD",x"FA",x"01",x"32",x"17",x"80", -- 0x0118
    x"3A",x"06",x"80",x"CD",x"F1",x"01",x"32",x"12", -- 0x0120
    x"80",x"3A",x"08",x"80",x"CD",x"F1",x"01",x"32", -- 0x0128
    x"13",x"80",x"3A",x"0A",x"80",x"CD",x"F1",x"01", -- 0x0130
    x"32",x"14",x"80",x"CD",x"FA",x"01",x"32",x"18", -- 0x0138
    x"80",x"B7",x"28",x"63",x"3A",x"17",x"80",x"B7", -- 0x0140
    x"28",x"79",x"3A",x"18",x"80",x"21",x"06",x"80", -- 0x0148
    x"CD",x"E3",x"01",x"CD",x"F1",x"01",x"47",x"3A", -- 0x0150
    x"17",x"80",x"21",x"00",x"80",x"CD",x"E3",x"01", -- 0x0158
    x"CD",x"F1",x"01",x"B8",x"F2",x"C3",x"01",x"18", -- 0x0160
    x"3E",x"FE",x"01",x"28",x"17",x"FE",x"02",x"28", -- 0x0168
    x"1A",x"FE",x"03",x"28",x"1D",x"FE",x"04",x"28", -- 0x0170
    x"20",x"FE",x"05",x"28",x"23",x"3A",x"1A",x"80", -- 0x0178
    x"32",x"0A",x"80",x"C9",x"3A",x"1A",x"80",x"32", -- 0x0180
    x"00",x"80",x"C9",x"3A",x"1A",x"80",x"32",x"02", -- 0x0188
    x"80",x"C9",x"3A",x"1A",x"80",x"32",x"04",x"80", -- 0x0190
    x"C9",x"3A",x"1A",x"80",x"32",x"06",x"80",x"C9", -- 0x0198
    x"3A",x"1A",x"80",x"32",x"08",x"80",x"C9",x"3A", -- 0x01A0
    x"17",x"80",x"B7",x"C8",x"FE",x"01",x"28",x"09", -- 0x01A8
    x"FE",x"02",x"28",x"0A",x"21",x"04",x"80",x"18", -- 0x01B0
    x"18",x"21",x"00",x"80",x"18",x"13",x"21",x"02", -- 0x01B8
    x"80",x"18",x"0E",x"3A",x"18",x"80",x"FE",x"01", -- 0x01C0
    x"28",x"0F",x"FE",x"02",x"28",x"10",x"21",x"0A", -- 0x01C8
    x"80",x"3A",x"1A",x"80",x"77",x"23",x"36",x"00", -- 0x01D0
    x"C9",x"21",x"06",x"80",x"18",x"F3",x"21",x"08", -- 0x01D8
    x"80",x"18",x"EE",x"FE",x"01",x"28",x"08",x"23", -- 0x01E0
    x"23",x"FE",x"02",x"28",x"02",x"23",x"23",x"7E", -- 0x01E8
    x"C9",x"21",x"42",x"02",x"5F",x"16",x"00",x"19", -- 0x01F0
    x"7E",x"C9",x"3A",x"12",x"80",x"21",x"13",x"80", -- 0x01F8
    x"BE",x"FA",x"15",x"02",x"3A",x"14",x"80",x"BE", -- 0x0200
    x"FA",x"34",x"02",x"3A",x"15",x"80",x"BE",x"FA", -- 0x0208
    x"40",x"02",x"3E",x"02",x"C9",x"21",x"14",x"80", -- 0x0210
    x"BE",x"FA",x"26",x"02",x"3A",x"15",x"80",x"BE", -- 0x0218
    x"FA",x"32",x"02",x"3E",x"03",x"C9",x"21",x"15", -- 0x0220
    x"80",x"BE",x"FA",x"2F",x"02",x"AF",x"C9",x"3E", -- 0x0228
    x"01",x"C9",x"AF",x"C9",x"21",x"15",x"80",x"BE", -- 0x0230
    x"FA",x"3D",x"02",x"AF",x"C9",x"3E",x"03",x"C9", -- 0x0238
    x"AF",x"C9",x"00",x"01",x"02",x"03",x"04",x"05", -- 0x0240
    x"06",x"07",x"08",x"09",x"0A",x"0B",x"0C",x"0D", -- 0x0248
    x"0E",x"0F",x"10",x"11",x"12",x"13",x"14",x"15", -- 0x0250
    x"16",x"17",x"18",x"19",x"1A",x"1B",x"1C",x"1D", -- 0x0258
    x"1E",x"1F",x"20",x"21",x"22",x"23",x"24",x"25", -- 0x0260
    x"26",x"27",x"28",x"29",x"2A",x"2B",x"2C",x"2D", -- 0x0268
    x"2E",x"2F",x"06",x"00",x"21",x"00",x"80",x"70", -- 0x0270
    x"23",x"7C",x"FE",x"84",x"20",x"F9",x"31",x"00", -- 0x0278
    x"84",x"ED",x"56",x"21",x"00",x"90",x"22",x"0C", -- 0x0280
    x"80",x"77",x"3E",x"07",x"D3",x"40",x"3E",x"3F", -- 0x0288
    x"32",x"0E",x"80",x"D3",x"80",x"3E",x"07",x"D3", -- 0x0290
    x"10",x"3E",x"3F",x"32",x"0F",x"80",x"D3",x"20", -- 0x0298
    x"CD",x"2D",x"04",x"CD",x"35",x"04",x"CD",x"3D", -- 0x02A0
    x"04",x"CD",x"45",x"04",x"CD",x"4D",x"04",x"CD", -- 0x02A8
    x"55",x"04",x"FB",x"3E",x"0F",x"D3",x"40",x"DB", -- 0x02B0
    x"80",x"E6",x"80",x"20",x"F6",x"3E",x"0F",x"D3", -- 0x02B8
    x"40",x"DB",x"80",x"E6",x"80",x"28",x"F6",x"F3", -- 0x02C0
    x"3E",x"01",x"32",x"10",x"80",x"3A",x"01",x"80", -- 0x02C8
    x"B7",x"CA",x"4B",x"03",x"3A",x"00",x"80",x"CD", -- 0x02D0
    x"04",x"08",x"FB",x"00",x"00",x"F3",x"3E",x"02", -- 0x02D8
    x"32",x"10",x"80",x"3A",x"03",x"80",x"B7",x"CA", -- 0x02E0
    x"54",x"03",x"3A",x"02",x"80",x"CD",x"04",x"08", -- 0x02E8
    x"FB",x"00",x"00",x"F3",x"3E",x"03",x"32",x"10", -- 0x02F0
    x"80",x"3A",x"05",x"80",x"B7",x"CA",x"5D",x"03", -- 0x02F8
    x"3A",x"04",x"80",x"CD",x"04",x"08",x"FB",x"00", -- 0x0300
    x"00",x"F3",x"3E",x"04",x"32",x"10",x"80",x"3A", -- 0x0308
    x"07",x"80",x"B7",x"CA",x"66",x"03",x"3A",x"06", -- 0x0310
    x"80",x"CD",x"04",x"08",x"FB",x"00",x"00",x"F3", -- 0x0318
    x"3E",x"05",x"32",x"10",x"80",x"3A",x"09",x"80", -- 0x0320
    x"B7",x"CA",x"6F",x"03",x"3A",x"08",x"80",x"CD", -- 0x0328
    x"04",x"08",x"FB",x"00",x"00",x"F3",x"3E",x"06", -- 0x0330
    x"32",x"10",x"80",x"3A",x"0B",x"80",x"B7",x"CA", -- 0x0338
    x"78",x"03",x"3A",x"0A",x"80",x"CD",x"04",x"08", -- 0x0340
    x"C3",x"B2",x"02",x"3A",x"00",x"80",x"CD",x"81", -- 0x0348
    x"03",x"C3",x"DA",x"02",x"3A",x"02",x"80",x"CD", -- 0x0350
    x"81",x"03",x"C3",x"F0",x"02",x"3A",x"04",x"80", -- 0x0358
    x"CD",x"81",x"03",x"C3",x"06",x"03",x"3A",x"06", -- 0x0360
    x"80",x"CD",x"81",x"03",x"C3",x"1C",x"03",x"3A", -- 0x0368
    x"08",x"80",x"CD",x"81",x"03",x"C3",x"32",x"03", -- 0x0370
    x"3A",x"0A",x"80",x"CD",x"81",x"03",x"C3",x"B2", -- 0x0378
    x"02",x"21",x"92",x"03",x"E5",x"87",x"5F",x"16", -- 0x0380
    x"00",x"21",x"CD",x"03",x"19",x"5E",x"23",x"56", -- 0x0388
    x"EB",x"E9",x"3A",x"10",x"80",x"FE",x"01",x"28", -- 0x0390
    x"16",x"FE",x"02",x"28",x"18",x"FE",x"03",x"28", -- 0x0398
    x"1A",x"FE",x"04",x"28",x"1C",x"FE",x"05",x"28", -- 0x03A0
    x"1E",x"3E",x"01",x"32",x"0B",x"80",x"C9",x"3E", -- 0x03A8
    x"01",x"32",x"01",x"80",x"C9",x"3E",x"01",x"32", -- 0x03B0
    x"03",x"80",x"C9",x"3E",x"01",x"32",x"05",x"80", -- 0x03B8
    x"C9",x"3E",x"01",x"32",x"07",x"80",x"C9",x"3E", -- 0x03C0
    x"01",x"32",x"09",x"80",x"C9",x"5D",x"04",x"C0", -- 0x03C8
    x"08",x"3C",x"09",x"B8",x"09",x"34",x"0A",x"B0", -- 0x03D0
    x"0A",x"F9",x"0C",x"1D",x"12",x"A9",x"13",x"B9", -- 0x03D8
    x"0D",x"C7",x"0D",x"2E",x"10",x"3C",x"10",x"43", -- 0x03E0
    x"10",x"B2",x"10",x"C0",x"10",x"00",x"00",x"00", -- 0x03E8
    x"00",x"00",x"11",x"3C",x"0B",x"E3",x"0B",x"6D", -- 0x03F0
    x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0400
    x"00",x"00",x"00",x"00",x"00",x"7A",x"0D",x"80", -- 0x0408
    x"11",x"19",x"12",x"B6",x"12",x"34",x"13",x"00", -- 0x0410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0418
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0420
    x"00",x"00",x"00",x"00",x"00",x"3E",x"08",x"D3", -- 0x0428
    x"40",x"AF",x"D3",x"80",x"C9",x"3E",x"09",x"D3", -- 0x0430
    x"40",x"AF",x"D3",x"80",x"C9",x"3E",x"0A",x"D3", -- 0x0438
    x"40",x"AF",x"D3",x"80",x"C9",x"3E",x"08",x"D3", -- 0x0440
    x"10",x"AF",x"D3",x"20",x"C9",x"3E",x"09",x"D3", -- 0x0448
    x"10",x"AF",x"D3",x"20",x"C9",x"3E",x"0A",x"D3", -- 0x0450
    x"10",x"AF",x"D3",x"20",x"C9",x"3A",x"10",x"80", -- 0x0458
    x"FE",x"01",x"28",x"19",x"FE",x"02",x"28",x"1E", -- 0x0460
    x"FE",x"03",x"28",x"23",x"FE",x"04",x"28",x"28", -- 0x0468
    x"FE",x"05",x"28",x"2D",x"06",x"24",x"CD",x"B8", -- 0x0470
    x"04",x"CD",x"55",x"04",x"C9",x"06",x"09",x"CD", -- 0x0478
    x"AA",x"04",x"CD",x"2D",x"04",x"C9",x"06",x"12", -- 0x0480
    x"CD",x"AA",x"04",x"CD",x"35",x"04",x"C9",x"06", -- 0x0488
    x"24",x"CD",x"AA",x"04",x"CD",x"3D",x"04",x"C9", -- 0x0490
    x"06",x"09",x"CD",x"B8",x"04",x"CD",x"45",x"04", -- 0x0498
    x"C9",x"06",x"12",x"CD",x"B8",x"04",x"CD",x"4D", -- 0x04A0
    x"04",x"C9",x"3E",x"07",x"D3",x"40",x"3A",x"0E", -- 0x04A8
    x"80",x"B0",x"32",x"0E",x"80",x"D3",x"80",x"C9", -- 0x04B0
    x"3E",x"07",x"D3",x"10",x"3A",x"0F",x"80",x"B0", -- 0x04B8
    x"32",x"0F",x"80",x"D3",x"20",x"C9",x"3A",x"10", -- 0x04C0
    x"80",x"FE",x"01",x"28",x"20",x"FE",x"02",x"28", -- 0x04C8
    x"2C",x"FE",x"03",x"28",x"2C",x"FE",x"04",x"28", -- 0x04D0
    x"2C",x"FE",x"05",x"28",x"2C",x"06",x"04",x"78", -- 0x04D8
    x"D3",x"10",x"7D",x"D3",x"20",x"04",x"78",x"D3", -- 0x04E0
    x"10",x"7C",x"D3",x"20",x"C9",x"06",x"00",x"78", -- 0x04E8
    x"D3",x"40",x"7D",x"D3",x"80",x"04",x"78",x"D3", -- 0x04F0
    x"40",x"7C",x"D3",x"80",x"C9",x"06",x"02",x"18", -- 0x04F8
    x"EE",x"06",x"04",x"18",x"EA",x"06",x"00",x"18", -- 0x0500
    x"D6",x"06",x"02",x"18",x"D2",x"3A",x"10",x"80", -- 0x0508
    x"FE",x"01",x"28",x"18",x"FE",x"02",x"28",x"1C", -- 0x0510
    x"FE",x"03",x"28",x"1E",x"FE",x"04",x"28",x"20", -- 0x0518
    x"FE",x"05",x"28",x"22",x"16",x"FB",x"1E",x"20", -- 0x0520
    x"CD",x"71",x"05",x"C9",x"16",x"FE",x"1E",x"08", -- 0x0528
    x"CD",x"62",x"05",x"C9",x"16",x"FD",x"1E",x"10", -- 0x0530
    x"18",x"F6",x"16",x"FB",x"1E",x"20",x"18",x"F0", -- 0x0538
    x"16",x"FE",x"1E",x"08",x"18",x"E2",x"16",x"FD", -- 0x0540
    x"1E",x"10",x"18",x"DC",x"3A",x"10",x"80",x"FE", -- 0x0548
    x"04",x"FA",x"5B",x"05",x"7A",x"D3",x"10",x"7B", -- 0x0550
    x"D3",x"20",x"C9",x"7A",x"D3",x"40",x"7B",x"D3", -- 0x0558
    x"80",x"C9",x"3E",x"07",x"D3",x"40",x"3A",x"0E", -- 0x0560
    x"80",x"A2",x"B3",x"32",x"0E",x"80",x"D3",x"80", -- 0x0568
    x"C9",x"3E",x"07",x"D3",x"10",x"3A",x"0F",x"80", -- 0x0570
    x"A2",x"B3",x"32",x"0F",x"80",x"D3",x"20",x"C9", -- 0x0578
    x"3A",x"10",x"80",x"FE",x"01",x"28",x"18",x"FE", -- 0x0580
    x"02",x"28",x"1C",x"FE",x"03",x"28",x"1E",x"FE", -- 0x0588
    x"04",x"28",x"20",x"FE",x"05",x"28",x"22",x"16", -- 0x0590
    x"DF",x"1E",x"04",x"CD",x"71",x"05",x"C9",x"16", -- 0x0598
    x"F7",x"1E",x"01",x"CD",x"62",x"05",x"C9",x"16", -- 0x05A0
    x"EF",x"1E",x"02",x"18",x"F6",x"16",x"DF",x"1E", -- 0x05A8
    x"04",x"18",x"F0",x"16",x"F7",x"1E",x"01",x"18", -- 0x05B0
    x"E2",x"16",x"EF",x"1E",x"02",x"18",x"DC",x"3A", -- 0x05B8
    x"10",x"80",x"FE",x"01",x"28",x"18",x"FE",x"02", -- 0x05C0
    x"28",x"1C",x"FE",x"03",x"28",x"1E",x"FE",x"04", -- 0x05C8
    x"28",x"20",x"FE",x"05",x"28",x"22",x"16",x"DB", -- 0x05D0
    x"1E",x"00",x"CD",x"71",x"05",x"C9",x"16",x"F6", -- 0x05D8
    x"1E",x"00",x"CD",x"62",x"05",x"C9",x"16",x"ED", -- 0x05E0
    x"1E",x"00",x"18",x"F6",x"16",x"DB",x"1E",x"00", -- 0x05E8
    x"18",x"F0",x"16",x"F6",x"1E",x"00",x"18",x"E2", -- 0x05F0
    x"16",x"ED",x"1E",x"00",x"18",x"DC",x"3A",x"10", -- 0x05F8
    x"80",x"FE",x"01",x"28",x"18",x"FE",x"02",x"28", -- 0x0600
    x"1C",x"FE",x"03",x"28",x"1C",x"FE",x"04",x"28", -- 0x0608
    x"1C",x"FE",x"05",x"28",x"1C",x"3E",x"0A",x"D3", -- 0x0610
    x"10",x"78",x"D3",x"20",x"C9",x"3E",x"08",x"D3", -- 0x0618
    x"40",x"78",x"D3",x"80",x"C9",x"3E",x"09",x"18", -- 0x0620
    x"F6",x"3E",x"0A",x"18",x"F2",x"3E",x"08",x"18", -- 0x0628
    x"E6",x"3E",x"09",x"18",x"E2",x"3A",x"10",x"80", -- 0x0630
    x"FE",x"04",x"FA",x"44",x"06",x"7A",x"D3",x"10", -- 0x0638
    x"DB",x"20",x"5F",x"C9",x"7A",x"D3",x"40",x"DB", -- 0x0640
    x"80",x"5F",x"C9",x"3A",x"10",x"80",x"FE",x"01", -- 0x0648
    x"28",x"17",x"FE",x"02",x"28",x"1A",x"FE",x"03", -- 0x0650
    x"28",x"1A",x"FE",x"04",x"28",x"1A",x"FE",x"05", -- 0x0658
    x"28",x"1A",x"3E",x"0A",x"D3",x"10",x"DB",x"20", -- 0x0660
    x"C9",x"3E",x"08",x"D3",x"40",x"DB",x"80",x"C9", -- 0x0668
    x"3E",x"09",x"18",x"F7",x"3E",x"0A",x"18",x"F3", -- 0x0670
    x"3E",x"08",x"18",x"E8",x"3E",x"09",x"18",x"E4", -- 0x0678
    x"3A",x"10",x"80",x"FE",x"01",x"28",x"20",x"FE", -- 0x0680
    x"02",x"28",x"2C",x"FE",x"03",x"28",x"2C",x"FE", -- 0x0688
    x"04",x"28",x"2C",x"FE",x"05",x"28",x"2C",x"06", -- 0x0690
    x"04",x"78",x"D3",x"10",x"DB",x"20",x"6F",x"04", -- 0x0698
    x"78",x"D3",x"10",x"DB",x"20",x"67",x"C9",x"06", -- 0x06A0
    x"00",x"78",x"D3",x"40",x"DB",x"80",x"6F",x"04", -- 0x06A8
    x"78",x"D3",x"40",x"DB",x"80",x"67",x"C9",x"06", -- 0x06B0
    x"02",x"18",x"EE",x"06",x"04",x"18",x"EA",x"06", -- 0x06B8
    x"00",x"18",x"D6",x"06",x"02",x"18",x"D2",x"3A", -- 0x06C0
    x"10",x"80",x"FE",x"04",x"28",x"21",x"FE",x"05", -- 0x06C8
    x"28",x"22",x"FE",x"06",x"28",x"23",x"FE",x"01", -- 0x06D0
    x"28",x"24",x"FE",x"02",x"28",x"25",x"11",x"FF", -- 0x06D8
    x"F3",x"2A",x"0C",x"80",x"7A",x"A4",x"67",x"7B", -- 0x06E0
    x"A5",x"6F",x"22",x"0C",x"80",x"77",x"C9",x"11", -- 0x06E8
    x"FC",x"FF",x"18",x"ED",x"11",x"F3",x"FF",x"18", -- 0x06F0
    x"E8",x"11",x"CF",x"FF",x"18",x"E3",x"11",x"3F", -- 0x06F8
    x"FF",x"18",x"DE",x"11",x"FF",x"FC",x"18",x"D9", -- 0x0700
    x"3A",x"10",x"80",x"FE",x"04",x"28",x"20",x"FE", -- 0x0708
    x"05",x"28",x"21",x"FE",x"06",x"28",x"22",x"FE", -- 0x0710
    x"01",x"28",x"23",x"FE",x"02",x"28",x"24",x"11", -- 0x0718
    x"FF",x"F3",x"2A",x"0C",x"80",x"7A",x"A4",x"67", -- 0x0720
    x"7B",x"A5",x"6F",x"22",x"0C",x"80",x"C9",x"11", -- 0x0728
    x"FC",x"FF",x"18",x"EE",x"11",x"F3",x"FF",x"18", -- 0x0730
    x"E9",x"11",x"CF",x"FF",x"18",x"E4",x"11",x"3F", -- 0x0738
    x"FF",x"18",x"DF",x"11",x"FF",x"FC",x"18",x"DA", -- 0x0740
    x"CD",x"08",x"07",x"3A",x"10",x"80",x"FE",x"04", -- 0x0748
    x"28",x"17",x"FE",x"05",x"28",x"18",x"FE",x"06", -- 0x0750
    x"28",x"19",x"FE",x"01",x"28",x"1A",x"FE",x"02", -- 0x0758
    x"28",x"1B",x"11",x"00",x"08",x"CD",x"F6",x"07", -- 0x0760
    x"C9",x"11",x"02",x"00",x"18",x"F7",x"11",x"08", -- 0x0768
    x"00",x"18",x"F2",x"11",x"20",x"00",x"18",x"ED", -- 0x0770
    x"11",x"80",x"00",x"18",x"E8",x"11",x"00",x"02", -- 0x0778
    x"18",x"E3",x"CD",x"08",x"07",x"3A",x"10",x"80", -- 0x0780
    x"FE",x"04",x"28",x"17",x"FE",x"05",x"28",x"18", -- 0x0788
    x"FE",x"06",x"28",x"19",x"FE",x"01",x"28",x"1A", -- 0x0790
    x"FE",x"02",x"28",x"1B",x"11",x"00",x"04",x"CD", -- 0x0798
    x"F6",x"07",x"C9",x"11",x"01",x"00",x"18",x"F7", -- 0x07A0
    x"11",x"04",x"00",x"18",x"F2",x"11",x"10",x"00", -- 0x07A8
    x"18",x"ED",x"11",x"40",x"00",x"18",x"E8",x"11", -- 0x07B0
    x"00",x"01",x"18",x"E3",x"CD",x"08",x"07",x"3A", -- 0x07B8
    x"10",x"80",x"FE",x"04",x"28",x"17",x"FE",x"05", -- 0x07C0
    x"28",x"18",x"FE",x"06",x"28",x"19",x"FE",x"01", -- 0x07C8
    x"28",x"1A",x"FE",x"02",x"28",x"1B",x"11",x"00", -- 0x07D0
    x"0C",x"CD",x"F6",x"07",x"C9",x"11",x"03",x"00", -- 0x07D8
    x"18",x"F7",x"11",x"0C",x"00",x"18",x"F2",x"11", -- 0x07E0
    x"30",x"00",x"18",x"ED",x"11",x"C0",x"00",x"18", -- 0x07E8
    x"E8",x"11",x"00",x"03",x"18",x"E3",x"2A",x"0C", -- 0x07F0
    x"80",x"7A",x"B4",x"67",x"7B",x"B5",x"6F",x"22"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
