library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.project_pkg.all;
use work.target_pkg.all;

package platform_pkg is

	--  
	-- PACE constants which *MUST* be defined
	--

	constant PACE_VIDEO_NUM_BITMAPS		    : natural := 1;
	constant PACE_VIDEO_NUM_TILEMAPS	    : natural := 1;
	constant PACE_VIDEO_NUM_SPRITES 	    : natural := 64;
	constant PACE_VIDEO_H_SIZE				    : integer := 256;
	constant PACE_VIDEO_V_SIZE				    : integer := 240;
	constant PACE_VIDEO_L_CROP            : integer := 0;
	constant PACE_VIDEO_R_CROP            : integer := PACE_VIDEO_L_CROP;
  constant PACE_VIDEO_PIPELINE_DELAY    : integer := 5;
	
	constant PACE_INPUTS_NUM_BYTES        : integer := 7;
	
	constant CLK0_FREQ_MHz		            : natural := 
    PACE_CLKIN0 * PACE_CLK0_MULTIPLY_BY / PACE_CLK0_DIVIDE_BY;

  --
	-- Platform-specific constants (optional)
	--

	-- this CLUT is for debug only
	-- the real machine has a bank of clut (palette) registers
	type clut_typ is array (0 to 31) of std_logic_vector(7 downto 0);

	-- clut entries for TENNIS in-game palette	
	--constant clut : clut_typ :=
	--(
	--	-- tile palette
	--	X"17", X"0F", X"30", X"19", X"17", X"0F", X"30", X"27", 
	--	X"17", X"21", X"30", X"02", X"17", X"0F", X"30", X"02", 
	--	-- sprite palette
	--	X"17", X"0F", X"27", X"21", X"17", X"07", X"27", X"20", 
	--	X"17", X"39", X"0F", X"17", X"17", X"07", X"36", X"2B"
	--);
	
	-- clut entries for WRECKING CREW in-game palette	
	--constant clut : clut_typ :=
	--(
	--	-- tile palette
	--	X"0F", X"1B", X"27", X"16", X"0F", X"1B", X"10", X"0F", 
	--	X"0F", X"1B", X"00", X"0F", X"0F", X"1B", X"30", X"02", 
	--	-- sprite palette
	--	X"0F", X"27", X"02", X"16", X"0F", X"02", X"16", X"27", 
	--	X"0F", X"36", X"02", X"17", X"0F", X"06", X"14", X"30"
	--);

	-- clut entries for SUPER MARIO BROS in-game palette	
	constant clut : clut_typ :=
	(
		-- tile palette
		X"22", X"29", X"1A", X"0F", X"0F", X"36", X"17", X"0F", 
		X"0F", X"30", X"21", X"0F", X"0F", X"27", X"17", X"0F", 
		-- sprite palette
		X"22", X"16", X"27", X"18", X"0F", X"1A", X"30", X"27", 
		X"0F", X"16", X"30", X"27", X"0F", X"0F", X"36", X"17"
	);

	-- Palette : Table of RGB entries	

	type pal_entry_typ is array (0 to 2) of std_logic_vector(5 downto 0);
	type pal_typ is array (0 to 63) of pal_entry_typ;

	constant pal : pal_typ :=
	(
		-- PAL palette taken from NINTENDULATOR emulator
		0 => (0=>"100000", 1=>"100000", 2=>"100000"),
		1 => (0=>"000000", 1=>"001111", 2=>"101001"),
		2 => (0=>"000000", 1=>"000100", 2=>"101100"),
		3 => (0=>"010001", 1=>"000000", 2=>"100101"),
		4 => (0=>"101000", 1=>"000000", 2=>"010111"),
		5 => (0=>"110001", 1=>"000000", 2=>"001010"),
		6 => (0=>"101110", 1=>"000001", 2=>"000000"),
		7 => (0=>"100011", 1=>"000101", 2=>"000000"),
		8 => (0=>"010111", 1=>"001011", 2=>"000000"),
		9 => (0=>"000100", 1=>"010001", 2=>"000000"),
		10 => (0=>"000001", 1=>"010010", 2=>"000000"),
		11 => (0=>"000000", 1=>"010001", 2=>"001011"),
		12 => (0=>"000000", 1=>"010000", 2=>"011001"),
		14 => (0=>"000001", 1=>"000001", 2=>"000001"),
		15 => (0=>"000001", 1=>"000001", 2=>"000001"),
		16 => (0=>"110001", 1=>"110001", 2=>"110001"),
		17 => (0=>"000000", 1=>"011101", 2=>"111111"),
		18 => (0=>"001000", 1=>"010101", 2=>"111111"),
		19 => (0=>"100000", 1=>"001101", 2=>"111110"),
		20 => (0=>"111010", 1=>"001011", 2=>"101101"),
		21 => (0=>"111111", 1=>"001010", 2=>"010100"),
		22 => (0=>"111111", 1=>"001000", 2=>"000000"),
		23 => (0=>"110101", 1=>"001100", 2=>"000000"),
		24 => (0=>"110001", 1=>"011000", 2=>"000000"),
		25 => (0=>"001101", 1=>"100000", 2=>"000000"),
		26 => (0=>"000001", 1=>"100011", 2=>"000000"),
		27 => (0=>"000000", 1=>"100010", 2=>"010101"),
		28 => (0=>"000000", 1=>"100110", 2=>"110011"),
		29 => (0=>"001000", 1=>"001000", 2=>"001000"),
		30 => (0=>"000010", 1=>"000010", 2=>"000010"),
		31 => (0=>"000010", 1=>"000010", 2=>"000010"),
		32 => (0=>"111111", 1=>"111111", 2=>"111111"),
		33 => (0=>"000011", 1=>"110101", 2=>"111111"),
		34 => (0=>"011010", 1=>"101000", 2=>"111111"),
		35 => (0=>"110101", 1=>"100000", 2=>"111111"),
		36 => (0=>"111111", 1=>"010001", 2=>"111100"),
		37 => (0=>"111111", 1=>"011000", 2=>"100010"),
		38 => (0=>"111111", 1=>"100010", 2=>"001100"),
		39 => (0=>"111111", 1=>"100111", 2=>"000100"),
		40 => (0=>"111110", 1=>"101111", 2=>"001000"),
		41 => (0=>"100111", 1=>"111000", 2=>"000011"),
		42 => (0=>"001010", 1=>"111100", 2=>"001101"),
		43 => (0=>"000011", 1=>"111100", 2=>"101001"),
		44 => (0=>"000001", 1=>"111110", 2=>"111111"),
		45 => (0=>"010111", 1=>"010111", 2=>"010111"),
		46 => (0=>"000011", 1=>"000011", 2=>"000011"),
		47 => (0=>"000011", 1=>"000011", 2=>"000011"),
		48 => (0=>"111111", 1=>"111111", 2=>"111111"),
		49 => (0=>"101001", 1=>"111111", 2=>"111111"),
		50 => (0=>"101100", 1=>"111011", 2=>"111111"),
		51 => (0=>"110110", 1=>"101010", 2=>"111010"),
		52 => (0=>"111111", 1=>"101010", 2=>"111110"),
		53 => (0=>"111111", 1=>"101010", 2=>"101100"),
		54 => (0=>"111111", 1=>"110100", 2=>"101100"),
		55 => (0=>"111111", 1=>"111011", 2=>"101001"),
		56 => (0=>"111111", 1=>"111101", 2=>"100111"),
		57 => (0=>"110101", 1=>"111010", 2=>"100101"),
		58 => (0=>"101001", 1=>"111011", 2=>"101011"),
		59 => (0=>"101000", 1=>"111100", 2=>"110110"),
		60 => (0=>"100110", 1=>"111111", 2=>"111111"),
		61 => (0=>"110111", 1=>"110111", 2=>"110111"),
		62 => (0=>"000100", 1=>"000100", 2=>"000100"),
		63 => (0=>"000100", 1=>"000100", 2=>"000100"),
		others => (others => (others => '0'))
	);

  type from_PLATFORM_IO_t is record
    not_used  : std_logic;
  end record;

  type to_PLATFORM_IO_t is record
    not_used  : std_logic;
  end record;

end;
