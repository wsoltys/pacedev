library work;
use work.pace_pkg.all;
use work.project_pkg.all;

package body platform_pkg is

  constant TUTANKHAM_SOURCE_ROOT_DIR  : string := "../../../../../src/platform/tutankhm/";

end platform_pkg;
