-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_PGM_01 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_PGM_01 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"AF",x"32",x"01",x"68",x"C3",x"D1",x"00",x"FF", -- 0x0000
    x"77",x"3C",x"23",x"77",x"3C",x"19",x"C9",x"FF", -- 0x0008
    x"77",x"23",x"10",x"FC",x"C9",x"FF",x"FF",x"FF", -- 0x0010
    x"77",x"23",x"10",x"FC",x"0D",x"20",x"F9",x"C9", -- 0x0018
    x"85",x"6F",x"3E",x"00",x"8C",x"67",x"7E",x"C9", -- 0x0020
    x"87",x"E1",x"5F",x"16",x"00",x"19",x"5E",x"23", -- 0x0028
    x"56",x"EB",x"E9",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0030
    x"E5",x"26",x"40",x"3A",x"A0",x"40",x"6F",x"CB", -- 0x0038
    x"7E",x"28",x"0E",x"72",x"2C",x"73",x"2C",x"7D", -- 0x0040
    x"FE",x"C0",x"30",x"02",x"3E",x"C0",x"32",x"A0", -- 0x0048
    x"40",x"E1",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C3",x"43", -- 0x0060
    x"0D",x"BC",x"4A",x"6E",x"40",x"40",x"53",x"54", -- 0x0068
    x"45",x"52",x"4E",x"40",x"40",x"31",x"39",x"38", -- 0x0070
    x"31",x"3F",x"BC",x"4A",x"6E",x"40",x"4B",x"4F", -- 0x0078
    x"4E",x"41",x"4D",x"49",x"40",x"40",x"31",x"39", -- 0x0080
    x"38",x"31",x"3F",x"54",x"4B",x"40",x"4F",x"55", -- 0x0088
    x"52",x"40",x"53",x"43",x"52",x"41",x"4D",x"42", -- 0x0090
    x"4C",x"45",x"40",x"53",x"59",x"53",x"54",x"45", -- 0x0098
    x"4D",x"40",x"02",x"3F",x"D5",x"4A",x"32",x"40", -- 0x00A0
    x"43",x"4F",x"49",x"4E",x"53",x"40",x"31",x"40", -- 0x00A8
    x"50",x"4C",x"41",x"59",x"3F",x"D5",x"4A",x"33", -- 0x00B0
    x"40",x"43",x"4F",x"49",x"4E",x"53",x"40",x"31", -- 0x00B8
    x"40",x"50",x"4C",x"41",x"59",x"3F",x"AF",x"01", -- 0x00C0
    x"02",x"04",x"32",x"02",x"82",x"81",x"10",x"FA", -- 0x00C8
    x"C9",x"3E",x"9B",x"32",x"03",x"81",x"3E",x"88", -- 0x00D0
    x"32",x"03",x"82",x"31",x"00",x"48",x"CD",x"C6", -- 0x00D8
    x"00",x"3A",x"02",x"81",x"17",x"38",x"F7",x"21", -- 0x00E0
    x"00",x"40",x"01",x"00",x"08",x"71",x"2C",x"20", -- 0x00E8
    x"FC",x"78",x"17",x"32",x"02",x"82",x"24",x"10", -- 0x00F0
    x"F4",x"3E",x"08",x"32",x"42",x"42",x"32",x"01", -- 0x00F8
    x"82",x"31",x"00",x"48",x"21",x"C0",x"40",x"06", -- 0x0100
    x"40",x"3E",x"FF",x"D7",x"21",x"43",x"42",x"06", -- 0x0108
    x"1C",x"D7",x"21",x"43",x"43",x"22",x"40",x"42", -- 0x0110
    x"3A",x"00",x"70",x"AF",x"32",x"01",x"68",x"32", -- 0x0118
    x"05",x"70",x"32",x"06",x"68",x"32",x"07",x"68", -- 0x0120
    x"32",x"02",x"82",x"21",x"C0",x"C0",x"22",x"A0", -- 0x0128
    x"40",x"3C",x"32",x"04",x"68",x"21",x"00",x"48", -- 0x0130
    x"22",x"0B",x"40",x"3E",x"20",x"32",x"08",x"40", -- 0x0138
    x"3E",x"10",x"32",x"17",x"40",x"3A",x"02",x"81", -- 0x0140
    x"0F",x"47",x"E6",x"03",x"32",x"00",x"40",x"78", -- 0x0148
    x"0F",x"0F",x"E6",x"01",x"32",x"0F",x"40",x"3A", -- 0x0150
    x"01",x"81",x"E6",x"03",x"FE",x"03",x"28",x"07", -- 0x0158
    x"C6",x"03",x"32",x"07",x"40",x"18",x"05",x"3E", -- 0x0160
    x"FF",x"32",x"07",x"40",x"CD",x"8E",x"30",x"AF", -- 0x0168
    x"3D",x"20",x"FD",x"CD",x"9D",x"30",x"06",x"04", -- 0x0170
    x"D9",x"CD",x"C6",x"00",x"D9",x"10",x"F9",x"3E", -- 0x0178
    x"28",x"07",x"C6",x"32",x"67",x"E6",x"0F",x"6F", -- 0x0180
    x"C6",x"63",x"77",x"01",x"02",x"0B",x"1E",x"09", -- 0x0188
    x"4F",x"57",x"70",x"06",x"03",x"DD",x"4E",x"03", -- 0x0190
    x"10",x"FB",x"77",x"59",x"06",x"FA",x"80",x"77", -- 0x0198
    x"0E",x"10",x"06",x"20",x"81",x"80",x"7E",x"FE", -- 0x01A0
    x"6F",x"C0",x"31",x"00",x"48",x"CD",x"C6",x"00", -- 0x01A8
    x"3A",x"02",x"81",x"17",x"30",x"F7",x"21",x"00", -- 0x01B0
    x"50",x"01",x"00",x"01",x"16",x"00",x"72",x"23", -- 0x01B8
    x"0B",x"78",x"B1",x"20",x"F9",x"16",x"3F",x"21", -- 0x01C0
    x"00",x"48",x"01",x"00",x"08",x"72",x"3A",x"00", -- 0x01C8
    x"70",x"23",x"0B",x"78",x"B1",x"20",x"F6",x"CD", -- 0x01D0
    x"03",x"02",x"30",x"22",x"CD",x"03",x"02",x"30", -- 0x01D8
    x"1D",x"3E",x"01",x"32",x"01",x"68",x"21",x"00", -- 0x01E0
    x"42",x"06",x"0A",x"36",x"00",x"2C",x"36",x"00", -- 0x01E8
    x"2C",x"36",x"01",x"2C",x"10",x"F5",x"21",x"AA", -- 0x01F0
    x"40",x"36",x"01",x"C3",x"17",x"02",x"3A",x"00", -- 0x01F8
    x"70",x"18",x"FB",x"0B",x"3A",x"00",x"70",x"3A", -- 0x0200
    x"01",x"81",x"07",x"D0",x"78",x"B1",x"20",x"F3", -- 0x0208
    x"3A",x"02",x"81",x"07",x"D0",x"37",x"C9",x"26", -- 0x0210
    x"40",x"3A",x"A1",x"40",x"6F",x"7E",x"87",x"30", -- 0x0218
    x"05",x"CD",x"5A",x"02",x"18",x"F1",x"E6",x"0F", -- 0x0220
    x"4F",x"06",x"00",x"36",x"FF",x"23",x"5E",x"36", -- 0x0228
    x"FF",x"2C",x"7D",x"FE",x"C0",x"30",x"02",x"3E", -- 0x0230
    x"C0",x"32",x"A1",x"40",x"7B",x"21",x"4A",x"02", -- 0x0238
    x"09",x"5E",x"23",x"56",x"21",x"17",x"02",x"E5", -- 0x0240
    x"EB",x"E9",x"C0",x"02",x"C1",x"02",x"C2",x"02", -- 0x0248
    x"20",x"03",x"B6",x"03",x"D2",x"03",x"19",x"04", -- 0x0250
    x"DE",x"06",x"3A",x"5F",x"42",x"47",x"E6",x"0F", -- 0x0258
    x"CA",x"79",x"02",x"21",x"19",x"40",x"CB",x"46", -- 0x0260
    x"C8",x"E6",x"03",x"CA",x"0C",x"0C",x"3D",x"CA", -- 0x0268
    x"D7",x"0B",x"3D",x"CA",x"1C",x"0B",x"C3",x"D7", -- 0x0270
    x"0B",x"11",x"E0",x"FF",x"21",x"E0",x"48",x"3A", -- 0x0278
    x"0E",x"40",x"A7",x"28",x"22",x"36",x"02",x"CD", -- 0x0280
    x"B1",x"02",x"21",x"40",x"4B",x"CD",x"AF",x"02", -- 0x0288
    x"3A",x"0D",x"40",x"A7",x"21",x"40",x"4B",x"28", -- 0x0290
    x"03",x"21",x"E0",x"48",x"CB",x"60",x"C8",x"3A", -- 0x0298
    x"06",x"40",x"0F",x"D0",x"C3",x"B8",x"02",x"21", -- 0x02A0
    x"E0",x"48",x"CD",x"B8",x"02",x"18",x"DB",x"36", -- 0x02A8
    x"01",x"19",x"36",x"25",x"19",x"36",x"20",x"C9", -- 0x02B0
    x"3E",x"10",x"77",x"19",x"77",x"19",x"77",x"C9", -- 0x02B8
    x"C9",x"C9",x"3E",x"1A",x"06",x"0B",x"F5",x"C5", -- 0x02C0
    x"CD",x"19",x"04",x"C1",x"F1",x"3C",x"10",x"F6", -- 0x02C8
    x"21",x"87",x"49",x"11",x"20",x"00",x"06",x"0A", -- 0x02D0
    x"DD",x"21",x"00",x"42",x"DD",x"7E",x"00",x"4F", -- 0x02D8
    x"E6",x"0F",x"77",x"19",x"79",x"0F",x"0F",x"0F", -- 0x02E0
    x"0F",x"E6",x"0F",x"77",x"19",x"DD",x"23",x"DD", -- 0x02E8
    x"7E",x"00",x"4F",x"E6",x"0F",x"77",x"19",x"79", -- 0x02F0
    x"0F",x"0F",x"0F",x"0F",x"E6",x"0F",x"77",x"19", -- 0x02F8
    x"DD",x"23",x"DD",x"7E",x"00",x"4F",x"E6",x"0F", -- 0x0300
    x"77",x"19",x"79",x"0F",x"0F",x"0F",x"0F",x"E6", -- 0x0308
    x"0F",x"28",x"01",x"77",x"11",x"62",x"FF",x"19", -- 0x0310
    x"11",x"20",x"00",x"DD",x"23",x"10",x"BD",x"C9", -- 0x0318
    x"4F",x"3A",x"06",x"40",x"0F",x"D0",x"79",x"A7", -- 0x0320
    x"28",x"48",x"4F",x"CD",x"7D",x"03",x"87",x"81", -- 0x0328
    x"4F",x"06",x"00",x"21",x"8C",x"03",x"09",x"A7", -- 0x0330
    x"06",x"03",x"1A",x"8E",x"27",x"12",x"13",x"23", -- 0x0338
    x"10",x"F8",x"D5",x"3A",x"0D",x"40",x"0F",x"30", -- 0x0340
    x"02",x"3E",x"01",x"CD",x"D2",x"03",x"D1",x"1B", -- 0x0348
    x"21",x"AA",x"40",x"06",x"03",x"1A",x"BE",x"D8", -- 0x0350
    x"20",x"05",x"1B",x"2B",x"10",x"F7",x"C9",x"CD", -- 0x0358
    x"7D",x"03",x"21",x"A8",x"40",x"06",x"03",x"1A", -- 0x0360
    x"77",x"13",x"23",x"10",x"FA",x"3E",x"02",x"C3", -- 0x0368
    x"D2",x"03",x"CD",x"7D",x"03",x"21",x"AB",x"40", -- 0x0370
    x"A7",x"06",x"03",x"18",x"BD",x"F5",x"3A",x"0D", -- 0x0378
    x"40",x"11",x"A2",x"40",x"0F",x"30",x"03",x"11", -- 0x0380
    x"A5",x"40",x"F1",x"C9",x"00",x"00",x"00",x"50", -- 0x0388
    x"00",x"00",x"00",x"01",x"00",x"50",x"01",x"00", -- 0x0390
    x"80",x"00",x"00",x"00",x"01",x"00",x"00",x"02", -- 0x0398
    x"00",x"00",x"03",x"00",x"00",x"01",x"00",x"00", -- 0x03A0
    x"02",x"00",x"80",x"00",x"00",x"00",x"02",x"00", -- 0x03A8
    x"10",x"00",x"00",x"00",x"08",x"00",x"F5",x"21", -- 0x03B0
    x"A2",x"40",x"A7",x"28",x"09",x"21",x"A5",x"40", -- 0x03B8
    x"3D",x"28",x"03",x"21",x"A8",x"40",x"36",x"00", -- 0x03C0
    x"23",x"36",x"00",x"23",x"36",x"00",x"F1",x"C3", -- 0x03C8
    x"D2",x"03",x"21",x"A4",x"40",x"DD",x"21",x"81", -- 0x03D0
    x"4B",x"A7",x"28",x"11",x"21",x"A7",x"40",x"DD", -- 0x03D8
    x"21",x"21",x"49",x"3D",x"28",x"07",x"21",x"AA", -- 0x03E0
    x"40",x"DD",x"21",x"41",x"4A",x"11",x"E0",x"FF", -- 0x03E8
    x"06",x"03",x"0E",x"04",x"7E",x"0F",x"0F",x"0F", -- 0x03F0
    x"0F",x"CD",x"04",x"04",x"7E",x"CD",x"04",x"04", -- 0x03F8
    x"2B",x"10",x"F1",x"C9",x"E6",x"0F",x"28",x"08", -- 0x0400
    x"0E",x"00",x"DD",x"77",x"00",x"DD",x"19",x"C9", -- 0x0408
    x"79",x"A7",x"28",x"F6",x"3E",x"10",x"0D",x"18", -- 0x0410
    x"F1",x"87",x"F5",x"21",x"86",x"04",x"E6",x"7F", -- 0x0418
    x"5F",x"16",x"00",x"19",x"5E",x"23",x"56",x"EB", -- 0x0420
    x"5E",x"23",x"56",x"23",x"EB",x"01",x"E0",x"FF", -- 0x0428
    x"F1",x"38",x"0E",x"FA",x"4B",x"04",x"1A",x"FE", -- 0x0430
    x"3F",x"C8",x"D6",x"30",x"77",x"13",x"09",x"18", -- 0x0438
    x"F5",x"1A",x"FE",x"3F",x"C8",x"36",x"10",x"13", -- 0x0440
    x"09",x"18",x"F6",x"22",x"B5",x"40",x"ED",x"53", -- 0x0448
    x"B3",x"40",x"EB",x"7B",x"E6",x"1F",x"47",x"87", -- 0x0450
    x"C6",x"20",x"6F",x"26",x"40",x"22",x"B1",x"40", -- 0x0458
    x"CB",x"3B",x"CB",x"3B",x"7A",x"E6",x"03",x"0F", -- 0x0460
    x"0F",x"B3",x"E6",x"F8",x"4F",x"21",x"00",x"48", -- 0x0468
    x"78",x"85",x"6F",x"11",x"20",x"00",x"43",x"36", -- 0x0470
    x"10",x"19",x"10",x"FB",x"2A",x"B1",x"40",x"71", -- 0x0478
    x"3E",x"01",x"32",x"B0",x"40",x"C9",x"D0",x"04", -- 0x0480
    x"DD",x"04",x"F1",x"04",x"FE",x"04",x"0B",x"05", -- 0x0488
    x"18",x"05",x"27",x"05",x"40",x"05",x"47",x"05", -- 0x0490
    x"59",x"05",x"75",x"05",x"91",x"05",x"98",x"05", -- 0x0498
    x"A7",x"05",x"69",x"00",x"69",x"00",x"7A",x"00", -- 0x04A0
    x"7A",x"00",x"8B",x"00",x"A4",x"00",x"B5",x"00", -- 0x04A8
    x"B9",x"05",x"CA",x"05",x"DB",x"05",x"E5",x"05", -- 0x04B0
    x"F7",x"05",x"0C",x"06",x"20",x"06",x"33",x"06", -- 0x04B8
    x"46",x"06",x"59",x"06",x"6C",x"06",x"7F",x"06", -- 0x04C0
    x"92",x"06",x"A5",x"06",x"B8",x"06",x"CB",x"06", -- 0x04C8
    x"96",x"4A",x"47",x"41",x"4D",x"45",x"40",x"40", -- 0x04D0
    x"4F",x"56",x"45",x"52",x"3F",x"F1",x"4A",x"50", -- 0x04D8
    x"55",x"53",x"48",x"40",x"53",x"54",x"41",x"52", -- 0x04E0
    x"54",x"40",x"42",x"55",x"54",x"54",x"4F",x"4E", -- 0x04E8
    x"3F",x"94",x"4A",x"50",x"4C",x"41",x"59",x"45", -- 0x04F0
    x"52",x"40",x"4F",x"4E",x"45",x"3F",x"94",x"4A", -- 0x04F8
    x"50",x"4C",x"41",x"59",x"45",x"52",x"40",x"54", -- 0x0500
    x"57",x"4F",x"3F",x"80",x"4A",x"48",x"49",x"47", -- 0x0508
    x"48",x"40",x"53",x"43",x"4F",x"52",x"45",x"3F", -- 0x0510
    x"9F",x"4B",x"40",x"43",x"52",x"45",x"44",x"49", -- 0x0518
    x"54",x"40",x"40",x"40",x"40",x"40",x"3F",x"51", -- 0x0520
    x"4B",x"48",x"4F",x"57",x"40",x"46",x"41",x"52", -- 0x0528
    x"40",x"43",x"41",x"4E",x"40",x"59",x"4F",x"55", -- 0x0530
    x"40",x"49",x"4E",x"56",x"41",x"44",x"45",x"3F", -- 0x0538
    x"5E",x"4B",x"46",x"55",x"45",x"4C",x"3F",x"CC", -- 0x0540
    x"4A",x"43",x"4F",x"4E",x"47",x"52",x"41",x"54", -- 0x0548
    x"55",x"4C",x"41",x"54",x"49",x"4F",x"4E",x"53", -- 0x0550
    x"3F",x"6E",x"4B",x"59",x"4F",x"55",x"40",x"43", -- 0x0558
    x"4F",x"4D",x"50",x"4C",x"45",x"54",x"45",x"44", -- 0x0560
    x"40",x"59",x"4F",x"55",x"52",x"40",x"44",x"55", -- 0x0568
    x"54",x"49",x"45",x"53",x"3F",x"70",x"4B",x"47", -- 0x0570
    x"4F",x"4F",x"44",x"40",x"4C",x"55",x"43",x"4B", -- 0x0578
    x"40",x"4E",x"45",x"58",x"54",x"40",x"54",x"49", -- 0x0580
    x"4D",x"45",x"40",x"41",x"47",x"41",x"49",x"4E", -- 0x0588
    x"3F",x"26",x"4A",x"50",x"4C",x"41",x"59",x"3F", -- 0x0590
    x"A9",x"4A",x"5B",x"40",x"53",x"43",x"52",x"41", -- 0x0598
    x"4D",x"42",x"4C",x"45",x"40",x"5B",x"3F",x"C7", -- 0x05A0
    x"4A",x"5B",x"40",x"53",x"43",x"4F",x"52",x"45", -- 0x05A8
    x"40",x"54",x"41",x"42",x"4C",x"45",x"40",x"5B", -- 0x05B0
    x"3F",x"D5",x"4A",x"31",x"40",x"43",x"4F",x"49", -- 0x05B8
    x"4E",x"40",x"40",x"32",x"40",x"50",x"4C",x"41", -- 0x05C0
    x"59",x"3F",x"78",x"4B",x"42",x"4F",x"4E",x"55", -- 0x05C8
    x"53",x"40",x"4A",x"45",x"54",x"40",x"40",x"46", -- 0x05D0
    x"4F",x"52",x"3F",x"58",x"49",x"30",x"30",x"30", -- 0x05D8
    x"40",x"50",x"54",x"53",x"3F",x"D4",x"4A",x"4F", -- 0x05E0
    x"4E",x"45",x"40",x"50",x"4C",x"41",x"59",x"45", -- 0x05E8
    x"52",x"40",x"4F",x"4E",x"4C",x"59",x"3F",x"F4", -- 0x05F0
    x"4A",x"4F",x"4E",x"45",x"40",x"4F",x"52",x"40", -- 0x05F8
    x"54",x"57",x"4F",x"40",x"50",x"4C",x"41",x"59", -- 0x0600
    x"45",x"52",x"53",x"3F",x"04",x"4B",x"5B",x"40", -- 0x0608
    x"53",x"43",x"4F",x"52",x"45",x"40",x"52",x"41", -- 0x0610
    x"4E",x"4B",x"49",x"4E",x"47",x"40",x"5B",x"3F", -- 0x0618
    x"E7",x"4A",x"31",x"53",x"54",x"40",x"40",x"40", -- 0x0620
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"50", -- 0x0628
    x"54",x"53",x"3F",x"E9",x"4A",x"32",x"4E",x"44", -- 0x0630
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0638
    x"40",x"40",x"50",x"54",x"53",x"3F",x"EB",x"4A", -- 0x0640
    x"33",x"52",x"44",x"40",x"40",x"40",x"40",x"40", -- 0x0648
    x"40",x"40",x"40",x"40",x"40",x"50",x"54",x"53", -- 0x0650
    x"3F",x"ED",x"4A",x"34",x"54",x"48",x"40",x"40", -- 0x0658
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0660
    x"50",x"54",x"53",x"3F",x"EF",x"4A",x"35",x"54", -- 0x0668
    x"48",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0670
    x"40",x"40",x"40",x"50",x"54",x"53",x"3F",x"F1", -- 0x0678
    x"4A",x"36",x"54",x"48",x"40",x"40",x"40",x"40", -- 0x0680
    x"40",x"40",x"40",x"40",x"40",x"40",x"50",x"54", -- 0x0688
    x"53",x"3F",x"F3",x"4A",x"37",x"54",x"48",x"40", -- 0x0690
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x0698
    x"40",x"50",x"54",x"53",x"3F",x"F5",x"4A",x"38", -- 0x06A0
    x"54",x"48",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x06A8
    x"40",x"40",x"40",x"40",x"50",x"54",x"53",x"3F", -- 0x06B0
    x"F7",x"4A",x"39",x"54",x"48",x"40",x"40",x"40", -- 0x06B8
    x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"50", -- 0x06C0
    x"54",x"53",x"3F",x"F9",x"4A",x"31",x"30",x"54", -- 0x06C8
    x"48",x"40",x"40",x"40",x"40",x"40",x"40",x"40", -- 0x06D0
    x"40",x"40",x"50",x"54",x"53",x"3F",x"A7",x"CA", -- 0x06D8
    x"AC",x"0C",x"3D",x"CA",x"DE",x"0A",x"3D",x"CA", -- 0x06E0
    x"CA",x"0C",x"C3",x"87",x"0C",x"60",x"D1",x"60", -- 0x06E8
    x"D1",x"00",x"00",x"60",x"D1",x"60",x"D1",x"00", -- 0x06F0
    x"00",x"60",x"D1",x"60",x"D1",x"00",x"00",x"60", -- 0x06F8
    x"D1",x"60",x"D1",x"00",x"00",x"70",x"D1",x"70", -- 0x0700
    x"D1",x"00",x"01",x"60",x"D1",x"60",x"D1",x"00", -- 0x0708
    x"01",x"60",x"D1",x"60",x"D1",x"00",x"00",x"78", -- 0x0710
    x"D1",x"78",x"D1",x"00",x"01",x"60",x"D1",x"60", -- 0x0718
    x"D1",x"00",x"01",x"48",x"D1",x"48",x"D1",x"00", -- 0x0720
    x"00",x"58",x"D1",x"58",x"D1",x"00",x"01",x"48", -- 0x0728
    x"D1",x"48",x"D1",x"00",x"00",x"58",x"D1",x"58", -- 0x0730
    x"D1",x"00",x"01",x"58",x"D1",x"58",x"D1",x"00", -- 0x0738
    x"01",x"68",x"D1",x"68",x"D1",x"00",x"01",x"68", -- 0x0740
    x"D1",x"68",x"D1",x"00",x"02",x"78",x"D1",x"78", -- 0x0748
    x"D1",x"00",x"01",x"78",x"D1",x"78",x"D1",x"00", -- 0x0750
    x"01",x"88",x"D1",x"88",x"D1",x"00",x"01",x"88", -- 0x0758
    x"D1",x"88",x"D1",x"00",x"02",x"98",x"D1",x"98", -- 0x0760
    x"D1",x"00",x"01",x"98",x"D1",x"98",x"D1",x"00", -- 0x0768
    x"01",x"90",x"D1",x"90",x"D1",x"00",x"04",x"90", -- 0x0770
    x"D1",x"90",x"D1",x"00",x"04",x"90",x"D1",x"90", -- 0x0778
    x"D1",x"00",x"01",x"90",x"D1",x"90",x"D1",x"00", -- 0x0780
    x"00",x"A0",x"D1",x"A0",x"D1",x"00",x"01",x"80", -- 0x0788
    x"D1",x"80",x"D1",x"00",x"00",x"90",x"D1",x"90", -- 0x0790
    x"D1",x"00",x"01",x"70",x"D1",x"70",x"D1",x"00", -- 0x0798
    x"00",x"80",x"D1",x"80",x"D1",x"00",x"01",x"60", -- 0x07A0
    x"D1",x"60",x"D1",x"00",x"00",x"70",x"D1",x"70", -- 0x07A8
    x"D1",x"00",x"01",x"50",x"D1",x"50",x"D1",x"00", -- 0x07B0
    x"00",x"60",x"D1",x"60",x"D1",x"00",x"01",x"50", -- 0x07B8
    x"D1",x"50",x"D1",x"00",x"00",x"48",x"D1",x"48", -- 0x07C0
    x"D1",x"00",x"00",x"58",x"D1",x"58",x"D1",x"00", -- 0x07C8
    x"01",x"50",x"D1",x"50",x"D1",x"00",x"00",x"50", -- 0x07D0
    x"D1",x"50",x"D1",x"00",x"00",x"60",x"D1",x"60", -- 0x07D8
    x"D1",x"00",x"01",x"58",x"D1",x"58",x"D1",x"00", -- 0x07E0
    x"00",x"68",x"D1",x"68",x"D1",x"00",x"01",x"60", -- 0x07E8
    x"D1",x"60",x"D1",x"00",x"00",x"70",x"D1",x"70", -- 0x07F0
    x"D1",x"00",x"01",x"68",x"D1",x"68",x"D1",x"00", -- 0x07F8
    x"00",x"78",x"D1",x"78",x"D1",x"00",x"01",x"70", -- 0x0800
    x"D1",x"70",x"D1",x"00",x"00",x"80",x"D1",x"80", -- 0x0808
    x"D1",x"00",x"01",x"80",x"D1",x"80",x"D1",x"00", -- 0x0810
    x"00",x"80",x"D1",x"80",x"D1",x"00",x"00",x"80", -- 0x0818
    x"D1",x"80",x"D1",x"00",x"04",x"80",x"D1",x"80", -- 0x0820
    x"D1",x"00",x"02",x"80",x"D1",x"80",x"D1",x"00", -- 0x0828
    x"04",x"80",x"D1",x"80",x"D1",x"00",x"01",x"80", -- 0x0830
    x"D1",x"80",x"D1",x"00",x"01",x"78",x"D1",x"78", -- 0x0838
    x"D1",x"00",x"01",x"70",x"D1",x"70",x"D1",x"00", -- 0x0840
    x"02",x"68",x"D1",x"68",x"D1",x"00",x"04",x"60", -- 0x0848
    x"D1",x"60",x"D1",x"00",x"01",x"60",x"D1",x"60", -- 0x0850
    x"D1",x"00",x"01",x"58",x"D1",x"58",x"D1",x"00", -- 0x0858
    x"00",x"58",x"D1",x"58",x"D1",x"00",x"00",x"60", -- 0x0860
    x"D1",x"60",x"D1",x"00",x"01",x"48",x"D1",x"48", -- 0x0868
    x"D1",x"00",x"00",x"48",x"D1",x"48",x"D1",x"00", -- 0x0870
    x"00",x"50",x"D1",x"50",x"D1",x"00",x"01",x"48", -- 0x0878
    x"D1",x"48",x"D1",x"00",x"01",x"58",x"D1",x"58", -- 0x0880
    x"D1",x"00",x"01",x"48",x"D1",x"48",x"D1",x"00", -- 0x0888
    x"00",x"50",x"D1",x"50",x"D1",x"00",x"01",x"48", -- 0x0890
    x"D1",x"48",x"D1",x"00",x"00",x"60",x"D1",x"60", -- 0x0898
    x"D1",x"00",x"01",x"50",x"D1",x"50",x"D1",x"00", -- 0x08A0
    x"02",x"40",x"D1",x"40",x"D1",x"00",x"00",x"60", -- 0x08A8
    x"D1",x"60",x"D1",x"00",x"01",x"40",x"D1",x"40", -- 0x08B0
    x"D1",x"00",x"00",x"60",x"D1",x"60",x"D1",x"00", -- 0x08B8
    x"01",x"40",x"D1",x"40",x"D1",x"00",x"00",x"50", -- 0x08C0
    x"D1",x"50",x"D1",x"00",x"01",x"40",x"D1",x"40", -- 0x08C8
    x"D1",x"00",x"00",x"50",x"D1",x"50",x"D1",x"00", -- 0x08D0
    x"01",x"60",x"D1",x"60",x"D1",x"00",x"00",x"60", -- 0x08D8
    x"D1",x"60",x"D1",x"00",x"02",x"60",x"D1",x"60", -- 0x08E0
    x"D1",x"00",x"00",x"60",x"D1",x"60",x"D1",x"00", -- 0x08E8
    x"02",x"60",x"D1",x"60",x"D1",x"00",x"00",x"60", -- 0x08F0
    x"D1",x"60",x"D1",x"00",x"02",x"70",x"D1",x"70", -- 0x08F8
    x"D1",x"00",x"01",x"60",x"D1",x"60",x"D1",x"00", -- 0x0900
    x"01",x"60",x"D1",x"60",x"D1",x"00",x"00",x"78", -- 0x0908
    x"D1",x"78",x"D1",x"00",x"01",x"60",x"D1",x"60", -- 0x0910
    x"D1",x"00",x"01",x"48",x"D1",x"48",x"D1",x"00", -- 0x0918
    x"00",x"58",x"D1",x"58",x"D1",x"00",x"01",x"48", -- 0x0920
    x"D1",x"48",x"D1",x"00",x"00",x"58",x"D1",x"58", -- 0x0928
    x"D1",x"00",x"01",x"58",x"D1",x"58",x"D1",x"00", -- 0x0930
    x"01",x"68",x"D1",x"68",x"D1",x"00",x"01",x"68", -- 0x0938
    x"D1",x"68",x"D1",x"00",x"02",x"78",x"D1",x"78", -- 0x0940
    x"D1",x"00",x"01",x"78",x"D1",x"78",x"D1",x"00", -- 0x0948
    x"01",x"88",x"D1",x"88",x"D1",x"00",x"01",x"88", -- 0x0950
    x"D1",x"88",x"D1",x"00",x"02",x"98",x"D1",x"98", -- 0x0958
    x"D1",x"00",x"01",x"98",x"D1",x"98",x"D1",x"00", -- 0x0960
    x"01",x"90",x"D1",x"90",x"D1",x"00",x"04",x"90", -- 0x0968
    x"D1",x"90",x"D1",x"00",x"04",x"90",x"D1",x"90", -- 0x0970
    x"D1",x"00",x"01",x"90",x"D1",x"90",x"D1",x"00", -- 0x0978
    x"00",x"A0",x"D1",x"A0",x"D1",x"00",x"01",x"80", -- 0x0980
    x"D1",x"80",x"D1",x"00",x"00",x"90",x"D1",x"90", -- 0x0988
    x"D1",x"00",x"01",x"70",x"D1",x"70",x"D1",x"00", -- 0x0990
    x"00",x"80",x"D1",x"80",x"D1",x"00",x"01",x"60", -- 0x0998
    x"D1",x"60",x"D1",x"00",x"00",x"70",x"D1",x"70", -- 0x09A0
    x"D1",x"00",x"01",x"50",x"D1",x"50",x"D1",x"00", -- 0x09A8
    x"00",x"60",x"D1",x"60",x"D1",x"00",x"01",x"50", -- 0x09B0
    x"D1",x"50",x"D1",x"00",x"00",x"48",x"D1",x"48", -- 0x09B8
    x"D1",x"00",x"00",x"58",x"D1",x"58",x"D1",x"00", -- 0x09C0
    x"01",x"50",x"D1",x"50",x"D1",x"00",x"00",x"50", -- 0x09C8
    x"D1",x"50",x"D1",x"00",x"00",x"60",x"D1",x"60", -- 0x09D0
    x"D1",x"00",x"01",x"58",x"D1",x"58",x"D1",x"00", -- 0x09D8
    x"00",x"68",x"D1",x"68",x"D1",x"00",x"01",x"60", -- 0x09E0
    x"D1",x"60",x"D1",x"00",x"00",x"70",x"D1",x"70", -- 0x09E8
    x"D1",x"00",x"01",x"68",x"D1",x"68",x"D1",x"00", -- 0x09F0
    x"00",x"78",x"D1",x"78",x"D1",x"00",x"01",x"70", -- 0x09F8
    x"D1",x"70",x"D1",x"00",x"00",x"80",x"D1",x"80", -- 0x0A00
    x"D1",x"00",x"01",x"80",x"D1",x"80",x"D1",x"00", -- 0x0A08
    x"00",x"80",x"D1",x"80",x"D1",x"00",x"00",x"80", -- 0x0A10
    x"D1",x"80",x"D1",x"00",x"04",x"80",x"D1",x"80", -- 0x0A18
    x"D1",x"00",x"02",x"80",x"D1",x"80",x"D1",x"00", -- 0x0A20
    x"04",x"80",x"D1",x"80",x"D1",x"00",x"01",x"80", -- 0x0A28
    x"D1",x"80",x"D1",x"00",x"01",x"78",x"D1",x"78", -- 0x0A30
    x"D1",x"00",x"01",x"70",x"D1",x"70",x"D1",x"00", -- 0x0A38
    x"02",x"68",x"D1",x"68",x"D1",x"00",x"04",x"60", -- 0x0A40
    x"D1",x"60",x"D1",x"00",x"01",x"60",x"D1",x"60", -- 0x0A48
    x"D1",x"00",x"01",x"58",x"D1",x"58",x"D1",x"00", -- 0x0A50
    x"00",x"58",x"D1",x"58",x"D1",x"00",x"00",x"60", -- 0x0A58
    x"D1",x"60",x"D1",x"00",x"01",x"48",x"D1",x"48", -- 0x0A60
    x"D1",x"00",x"00",x"48",x"D1",x"48",x"D1",x"00", -- 0x0A68
    x"00",x"50",x"D1",x"50",x"D1",x"00",x"01",x"48", -- 0x0A70
    x"D1",x"48",x"D1",x"00",x"01",x"58",x"D1",x"58", -- 0x0A78
    x"D1",x"00",x"01",x"48",x"D1",x"48",x"D1",x"00", -- 0x0A80
    x"00",x"50",x"D1",x"50",x"D1",x"00",x"01",x"48", -- 0x0A88
    x"D1",x"48",x"D1",x"00",x"00",x"60",x"D1",x"60", -- 0x0A90
    x"D1",x"00",x"01",x"50",x"D1",x"50",x"D1",x"00", -- 0x0A98
    x"02",x"40",x"D1",x"40",x"D1",x"00",x"00",x"60", -- 0x0AA0
    x"D1",x"60",x"D1",x"00",x"01",x"40",x"D1",x"40", -- 0x0AA8
    x"D1",x"00",x"00",x"60",x"D1",x"60",x"D1",x"00", -- 0x0AB0
    x"01",x"40",x"D1",x"40",x"D1",x"00",x"00",x"50", -- 0x0AB8
    x"D1",x"50",x"D1",x"00",x"01",x"60",x"D1",x"60", -- 0x0AC0
    x"D1",x"00",x"00",x"60",x"D1",x"60",x"D1",x"00", -- 0x0AC8
    x"00",x"60",x"D1",x"60",x"D1",x"00",x"00",x"60", -- 0x0AD0
    x"D1",x"60",x"D1",x"00",x"00",x"FF",x"3E",x"05", -- 0x0AD8
    x"CD",x"19",x"04",x"3A",x"02",x"40",x"FE",x"63", -- 0x0AE0
    x"38",x"02",x"3E",x"63",x"CD",x"02",x"0B",x"47", -- 0x0AE8
    x"E6",x"F0",x"28",x"07",x"0F",x"0F",x"0F",x"0F", -- 0x0AF0
    x"32",x"9F",x"4A",x"78",x"E6",x"0F",x"32",x"7F", -- 0x0AF8
    x"4A",x"C9",x"47",x"E6",x"0F",x"C6",x"00",x"27", -- 0x0B00
    x"4F",x"78",x"E6",x"F0",x"28",x"0B",x"0F",x"0F", -- 0x0B08
    x"0F",x"0F",x"47",x"AF",x"C6",x"16",x"27",x"10", -- 0x0B10
    x"FB",x"81",x"27",x"C9",x"3A",x"10",x"41",x"0F", -- 0x0B18
    x"D0",x"3A",x"30",x"42",x"0F",x"D0",x"2A",x"35", -- 0x0B20
    x"42",x"7D",x"E6",x"E0",x"6F",x"11",x"05",x"00", -- 0x0B28
    x"19",x"3E",x"10",x"06",x"19",x"D7",x"11",x"07", -- 0x0B30
    x"00",x"19",x"06",x"19",x"D7",x"DD",x"21",x"30", -- 0x0B38
    x"42",x"DD",x"7E",x"01",x"DD",x"6E",x"02",x"DD", -- 0x0B40
    x"66",x"03",x"77",x"7D",x"E6",x"1F",x"47",x"3E", -- 0x0B48
    x"1D",x"90",x"28",x"10",x"47",x"0E",x"39",x"3A", -- 0x0B50
    x"1D",x"41",x"E6",x"1C",x"28",x"02",x"0E",x"3D", -- 0x0B58
    x"23",x"71",x"10",x"FC",x"DD",x"7E",x"04",x"DD", -- 0x0B60
    x"6E",x"05",x"DD",x"66",x"06",x"77",x"7D",x"E6", -- 0x0B68
    x"1F",x"47",x"3E",x"1D",x"90",x"28",x"10",x"47", -- 0x0B70
    x"0E",x"39",x"3A",x"1D",x"41",x"E6",x"1C",x"28", -- 0x0B78
    x"02",x"0E",x"D0",x"23",x"71",x"10",x"FC",x"DD", -- 0x0B80
    x"36",x"00",x"00",x"DD",x"CB",x"08",x"46",x"C8", -- 0x0B88
    x"DD",x"7E",x"09",x"DD",x"6E",x"0A",x"DD",x"66", -- 0x0B90
    x"0B",x"77",x"7D",x"E6",x"1F",x"D6",x"05",x"28", -- 0x0B98
    x"10",x"47",x"0E",x"39",x"3A",x"1D",x"41",x"E6", -- 0x0BA0
    x"1C",x"28",x"02",x"0E",x"D0",x"2B",x"71",x"10", -- 0x0BA8
    x"FC",x"DD",x"7E",x"0C",x"DD",x"6E",x"0D",x"DD", -- 0x0BB0
    x"66",x"0E",x"77",x"7D",x"E6",x"1F",x"D6",x"05", -- 0x0BB8
    x"28",x"10",x"47",x"0E",x"39",x"3A",x"1D",x"41", -- 0x0BC0
    x"E6",x"1C",x"28",x"02",x"0E",x"3D",x"2B",x"71", -- 0x0BC8
    x"10",x"FC",x"DD",x"36",x"08",x"00",x"C9",x"11", -- 0x0BD0
    x"04",x"00",x"06",x"08",x"DD",x"21",x"60",x"42", -- 0x0BD8
    x"D9",x"CD",x"EA",x"0B",x"D9",x"DD",x"19",x"10", -- 0x0BE0
    x"F7",x"C9",x"DD",x"CB",x"00",x"46",x"C8",x"DD", -- 0x0BE8
    x"7E",x"01",x"87",x"87",x"DD",x"6E",x"02",x"DD", -- 0x0BF0
    x"66",x"03",x"77",x"3C",x"23",x"77",x"3C",x"11", -- 0x0BF8
    x"1F",x"00",x"19",x"77",x"3C",x"23",x"77",x"DD", -- 0x0C00
    x"36",x"00",x"00",x"C9",x"3A",x"05",x"41",x"0F", -- 0x0C08
    x"4F",x"E6",x"78",x"0F",x"0F",x"0F",x"47",x"3E", -- 0x0C10
    x"0F",x"90",x"21",x"BE",x"4A",x"11",x"E0",x"FF", -- 0x0C18
    x"04",x"05",x"28",x"05",x"36",x"CB",x"19",x"10", -- 0x0C20
    x"FB",x"47",x"79",x"E6",x"07",x"D9",x"21",x"41", -- 0x0C28
    x"0C",x"5F",x"16",x"00",x"19",x"7E",x"D9",x"77", -- 0x0C30
    x"04",x"05",x"C8",x"19",x"36",x"3C",x"10",x"FB", -- 0x0C38
    x"C9",x"3C",x"C4",x"C5",x"C6",x"C7",x"C8",x"C9", -- 0x0C40
    x"CA",x"CD",x"0C",x"0C",x"3A",x"01",x"41",x"21", -- 0x0C48
    x"64",x"4B",x"11",x"E0",x"FF",x"47",x"3E",x"18", -- 0x0C50
    x"90",x"04",x"05",x"28",x"05",x"36",x"0C",x"19", -- 0x0C58
    x"10",x"FB",x"47",x"A7",x"28",x"05",x"36",x"10", -- 0x0C60
    x"19",x"10",x"FB",x"3A",x"02",x"41",x"21",x"63", -- 0x0C68
    x"4B",x"47",x"3E",x"18",x"90",x"04",x"05",x"28", -- 0x0C70
    x"05",x"36",x"0D",x"19",x"10",x"FB",x"47",x"A7", -- 0x0C78
    x"C8",x"36",x"10",x"19",x"10",x"FB",x"C9",x"21", -- 0x0C80
    x"BF",x"4B",x"11",x"E0",x"FF",x"06",x"0C",x"36", -- 0x0C88
    x"10",x"19",x"10",x"FB",x"21",x"BF",x"4B",x"3A", -- 0x0C90
    x"08",x"41",x"A7",x"C8",x"FE",x"07",x"38",x"02", -- 0x0C98
    x"3E",x"06",x"47",x"36",x"0A",x"19",x"36",x"0B", -- 0x0CA0
    x"19",x"10",x"F8",x"C9",x"3A",x"00",x"41",x"E6", -- 0x0CA8
    x"0F",x"3C",x"47",x"3E",x"10",x"90",x"21",x"5F", -- 0x0CB0
    x"48",x"11",x"20",x"00",x"36",x"0E",x"19",x"10", -- 0x0CB8
    x"FB",x"A7",x"C8",x"36",x"10",x"19",x"3D",x"20", -- 0x0CC0
    x"FA",x"C9",x"DD",x"21",x"63",x"4B",x"11",x"E0", -- 0x0CC8
    x"FF",x"21",x"0B",x"0D",x"06",x"18",x"7E",x"DD", -- 0x0CD0
    x"77",x"00",x"23",x"DD",x"19",x"10",x"F7",x"21", -- 0x0CD8
    x"64",x"4B",x"11",x"E0",x"FF",x"DD",x"21",x"23", -- 0x0CE0
    x"0D",x"06",x"18",x"DD",x"7E",x"00",x"77",x"DD", -- 0x0CE8
    x"23",x"19",x"10",x"F7",x"3A",x"1E",x"41",x"3C", -- 0x0CF0
    x"47",x"21",x"64",x"4B",x"36",x"81",x"19",x"36", -- 0x0CF8
    x"82",x"19",x"36",x"82",x"19",x"36",x"83",x"19", -- 0x0D00
    x"10",x"F2",x"C9",x"50",x"51",x"52",x"6D",x"53", -- 0x0D08
    x"54",x"55",x"6D",x"56",x"57",x"55",x"6D",x"58", -- 0x0D10
    x"59",x"5A",x"6D",x"5B",x"59",x"5A",x"6D",x"64", -- 0x0D18
    x"65",x"51",x"66",x"6E",x"6F",x"6F",x"80",x"6E", -- 0x0D20
    x"6F",x"6F",x"80",x"6E",x"6F",x"6F",x"80",x"6E", -- 0x0D28
    x"6F",x"6F",x"80",x"6E",x"6F",x"6F",x"80",x"6E", -- 0x0D30
    x"6F",x"6F",x"80",x"6E",x"6F",x"6F",x"80",x"6E", -- 0x0D38
    x"6F",x"6F",x"80",x"F5",x"C5",x"D5",x"E5",x"08", -- 0x0D40
    x"D9",x"F5",x"C5",x"D5",x"E5",x"DD",x"E5",x"FD", -- 0x0D48
    x"E5",x"AF",x"32",x"01",x"68",x"21",x"20",x"40", -- 0x0D50
    x"11",x"00",x"50",x"01",x"80",x"00",x"ED",x"B0", -- 0x0D58
    x"3A",x"00",x"70",x"3A",x"15",x"40",x"32",x"16", -- 0x0D60
    x"40",x"3A",x"13",x"40",x"32",x"15",x"40",x"2A", -- 0x0D68
    x"10",x"40",x"22",x"13",x"40",x"21",x"12",x"40", -- 0x0D70
    x"3A",x"02",x"81",x"2F",x"77",x"2B",x"3A",x"01", -- 0x0D78
    x"81",x"2F",x"77",x"2B",x"3A",x"00",x"81",x"2F", -- 0x0D80
    x"77",x"21",x"5F",x"42",x"35",x"CD",x"B9",x"0D", -- 0x0D88
    x"CD",x"50",x"30",x"21",x"A5",x"0D",x"E5",x"3A", -- 0x0D90
    x"05",x"40",x"EF",x"7C",x"0E",x"7D",x"0F",x"B7", -- 0x0D98
    x"11",x"DE",x"12",x"F6",x"12",x"FD",x"E1",x"DD", -- 0x0DA0
    x"E1",x"E1",x"D1",x"C1",x"F1",x"D9",x"08",x"E1", -- 0x0DA8
    x"D1",x"C1",x"3E",x"01",x"32",x"01",x"68",x"F1", -- 0x0DB0
    x"C9",x"21",x"18",x"40",x"7E",x"A7",x"28",x"03", -- 0x0DB8
    x"35",x"3E",x"01",x"32",x"02",x"68",x"21",x"10", -- 0x0DC0
    x"40",x"7E",x"2C",x"2C",x"2C",x"B6",x"2C",x"2C", -- 0x0DC8
    x"2F",x"A6",x"2C",x"E6",x"C4",x"28",x"21",x"47", -- 0x0DD0
    x"E6",x"C0",x"28",x"05",x"3E",x"06",x"32",x"18", -- 0x0DD8
    x"40",x"CD",x"34",x"0E",x"21",x"02",x"40",x"7E", -- 0x0DE0
    x"FE",x"63",x"38",x"02",x"36",x"63",x"3A",x"06", -- 0x0DE8
    x"40",x"0F",x"38",x"04",x"11",x"01",x"07",x"FF", -- 0x0DF0
    x"21",x"03",x"40",x"5E",x"16",x"06",x"1A",x"1C", -- 0x0DF8
    x"73",x"23",x"86",x"3D",x"77",x"3A",x"B0",x"40", -- 0x0E00
    x"0F",x"D0",x"2A",x"B1",x"40",x"7E",x"E6",x"07", -- 0x0E08
    x"20",x"1B",x"EB",x"2A",x"B3",x"40",x"7E",x"FE", -- 0x0E10
    x"3F",x"28",x"11",x"23",x"22",x"B3",x"40",x"D6", -- 0x0E18
    x"30",x"2A",x"B5",x"40",x"77",x"01",x"E0",x"FF", -- 0x0E20
    x"09",x"22",x"B5",x"40",x"EB",x"35",x"C0",x"AF", -- 0x0E28
    x"32",x"B0",x"40",x"C9",x"3A",x"02",x"82",x"CB", -- 0x0E30
    x"67",x"28",x"03",x"E6",x"0F",x"C0",x"21",x"02", -- 0x0E38
    x"40",x"78",x"E6",x"84",x"28",x"0E",x"34",x"3A", -- 0x0E40
    x"00",x"40",x"A7",x"C8",x"34",x"3D",x"C8",x"34", -- 0x0E48
    x"3D",x"C8",x"34",x"C9",x"3A",x"00",x"40",x"2D", -- 0x0E50
    x"34",x"A7",x"28",x"08",x"3D",x"28",x"0A",x"3D", -- 0x0E58
    x"28",x"0C",x"18",x"0F",x"7E",x"FE",x"02",x"18", -- 0x0E60
    x"0D",x"7E",x"FE",x"01",x"18",x"08",x"7E",x"FE", -- 0x0E68
    x"03",x"18",x"03",x"7E",x"FE",x"04",x"D8",x"36", -- 0x0E70
    x"00",x"2C",x"34",x"C9",x"2A",x"0B",x"40",x"06", -- 0x0E78
    x"20",x"3E",x"10",x"D7",x"22",x"0B",x"40",x"21", -- 0x0E80
    x"08",x"40",x"35",x"C0",x"2D",x"2D",x"36",x"00", -- 0x0E88
    x"2D",x"36",x"01",x"AF",x"32",x"0A",x"40",x"21", -- 0x0E90
    x"BD",x"0E",x"CD",x"AD",x"0E",x"11",x"04",x"06", -- 0x0E98
    x"FF",x"11",x"00",x"05",x"FF",x"1E",x"02",x"FF", -- 0x0EA0
    x"AF",x"32",x"14",x"45",x"C9",x"11",x"20",x"40", -- 0x0EA8
    x"06",x"20",x"EB",x"36",x"00",x"2C",x"1A",x"77", -- 0x0EB0
    x"2C",x"13",x"10",x"F7",x"C9",x"00",x"05",x"00", -- 0x0EB8
    x"07",x"07",x"01",x"06",x"00",x"00",x"00",x"00", -- 0x0EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0ED0
    x"00",x"00",x"00",x"01",x"06",x"00",x"05",x"00", -- 0x0ED8
    x"00",x"01",x"01",x"06",x"03",x"03",x"04",x"04", -- 0x0EE0
    x"04",x"04",x"00",x"00",x"00",x"02",x"02",x"02", -- 0x0EE8
    x"00",x"00",x"00",x"04",x"04",x"04",x"04",x"04", -- 0x0EF0
    x"06",x"06",x"06",x"06",x"06",x"00",x"05",x"02", -- 0x0EF8
    x"02",x"02",x"02",x"02",x"06",x"06",x"06",x"06", -- 0x0F00
    x"06",x"06",x"06",x"06",x"06",x"04",x"04",x"04", -- 0x0F08
    x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"06", -- 0x0F10
    x"06",x"00",x"06",x"06",x"06",x"00",x"05",x"06", -- 0x0F18
    x"06",x"06",x"06",x"06",x"02",x"00",x"00",x"00", -- 0x0F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F30
    x"00",x"00",x"06",x"06",x"06",x"00",x"05",x"04", -- 0x0F38
    x"04",x"04",x"04",x"04",x"02",x"02",x"02",x"02", -- 0x0F40
    x"02",x"02",x"06",x"06",x"06",x"06",x"06",x"06", -- 0x0F48
    x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07", -- 0x0F50
    x"06",x"06",x"06",x"06",x"06",x"00",x"05",x"01", -- 0x0F58
    x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"03", -- 0x0F60
    x"03",x"04",x"04",x"05",x"05",x"06",x"06",x"07", -- 0x0F68
    x"07",x"01",x"01",x"02",x"02",x"01",x"01",x"01", -- 0x0F70
    x"01",x"01",x"01",x"01",x"06",x"21",x"A9",x"11", -- 0x0F78
    x"E5",x"3A",x"41",x"45",x"EF",x"99",x"0F",x"C7", -- 0x0F80
    x"0F",x"07",x"10",x"29",x"10",x"3E",x"10",x"DB", -- 0x0F88
    x"10",x"04",x"11",x"25",x"11",x"40",x"11",x"8C", -- 0x0F90
    x"11",x"3E",x"01",x"32",x"04",x"68",x"3D",x"32", -- 0x0F98
    x"03",x"68",x"AF",x"32",x"19",x"40",x"21",x"20", -- 0x0FA0
    x"40",x"11",x"21",x"40",x"01",x"7F",x"00",x"36", -- 0x0FA8
    x"00",x"ED",x"B0",x"21",x"02",x"48",x"22",x"0B", -- 0x0FB0
    x"40",x"21",x"09",x"40",x"36",x"20",x"21",x"41", -- 0x0FB8
    x"45",x"34",x"AF",x"32",x"06",x"40",x"C9",x"2A", -- 0x0FC0
    x"0B",x"40",x"06",x"1E",x"3E",x"10",x"D7",x"11", -- 0x0FC8
    x"02",x"00",x"19",x"22",x"0B",x"40",x"21",x"09", -- 0x0FD0
    x"40",x"35",x"C0",x"21",x"FD",x"0E",x"CD",x"AD", -- 0x0FD8
    x"0E",x"AF",x"32",x"06",x"68",x"32",x"07",x"68", -- 0x0FE0
    x"21",x"41",x"45",x"34",x"2D",x"36",x"00",x"11", -- 0x0FE8
    x"01",x"07",x"FF",x"11",x"06",x"06",x"FF",x"11", -- 0x0FF0
    x"12",x"06",x"FF",x"11",x"0F",x"06",x"FF",x"11"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
