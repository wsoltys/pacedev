library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

library work;
use work.pace_pkg.all;
use work.kbd_pkg.all;

entity inputmapper is
	generic
	(
			NUM_INPUTS	: positive := 2
	);
	port
	(
	    clk       : in std_logic;
	    rst_n     : in std_logic;

	    -- inputs from keyboard controller
	    reset     : in std_logic;
	    press     : in std_logic;
	    release   : in std_logic;
	    data      : in std_logic_vector(7 downto 0);
			-- inputs from jamma interface
			jamma			: in JAMMAInputsType;

	    -- user outputs
			dips			: in	std_logic_vector(7 downto 0);
			inputs		: out	in8(0 to NUM_INPUTS-1)
	);
end inputmapper;

architecture SYN of inputmapper is

begin

    latchInputs: process (clk, rst_n)

    begin

         -- note: all inputs are active LOW

        if rst_n = '0' then
					inputs(0) <= "10101111";
					inputs(1) <= (others => '1');
					inputs(2) <= (others => '1');
        elsif rising_edge (clk) then
          if (press or release) = '1' then
               case data(7 downto 0) is
                    -- IN0
										-- bit6 is vblank
                    when SCANCODE_S =>
                         inputs(0)(5) <= release;

                    -- IN1
                    when SCANCODE_5 =>
                         inputs(1)(7) <= release;
                    when SCANCODE_6 =>
                         inputs(1)(6) <= release;
                    when SCANCODE_7 =>
                         inputs(1)(5) <= release;
                    when SCANCODE_LCTRL =>
                         inputs(1)(2) <= release;
                    when SCANCODE_2 =>
                         inputs(1)(1) <= release;
                    when SCANCODE_1 =>
                         inputs(1)(0) <= release;

                    when others =>
               end case;
            end if; -- press or release
            if (reset = '1') then
							inputs(0) <= "10101111";
							inputs(1) <= (others => '1');
							inputs(2) <= (others => '1');
            end if;
        end if; -- rising_edge (clk)
    end process latchInputs;

end SYN;


