-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_OBJ_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_OBJ_0 is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"38",x"7C",x"C1",x"81",x"85",x"7C",x"38",x"00", -- 0x0000
    x"01",x"01",x"FD",x"FD",x"41",x"01",x"00",x"00", -- 0x0008
    x"61",x"F1",x"B9",x"99",x"9D",x"CD",x"45",x"00", -- 0x0010
    x"8C",x"DD",x"F1",x"B1",x"91",x"85",x"04",x"00", -- 0x0018
    x"08",x"FD",x"FD",x"C8",x"68",x"38",x"18",x"00", -- 0x0020
    x"1C",x"BD",x"A1",x"A1",x"A1",x"E5",x"E4",x"00", -- 0x0028
    x"0C",x"9D",x"91",x"91",x"D1",x"7D",x"3C",x"00", -- 0x0030
    x"C0",x"E0",x"B0",x"9D",x"8D",x"C0",x"C0",x"00", -- 0x0038
    x"0C",x"6D",x"99",x"99",x"B1",x"F1",x"6C",x"00", -- 0x0040
    x"78",x"FC",x"95",x"91",x"91",x"F1",x"60",x"00", -- 0x0048
    x"3D",x"7D",x"C8",x"88",x"C8",x"7D",x"3D",x"00", -- 0x0050
    x"6C",x"FD",x"91",x"91",x"91",x"FD",x"FD",x"00", -- 0x0058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0060
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00", -- 0x0068
    x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x0070
    x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0080
    x"3D",x"7D",x"C8",x"88",x"C8",x"7D",x"3D",x"00", -- 0x0088
    x"6C",x"FD",x"91",x"91",x"91",x"FD",x"FD",x"00", -- 0x0090
    x"44",x"C5",x"81",x"81",x"C5",x"7C",x"38",x"00", -- 0x0098
    x"38",x"7C",x"C5",x"81",x"81",x"FD",x"FD",x"00", -- 0x00A0
    x"81",x"91",x"91",x"91",x"FD",x"FD",x"00",x"00", -- 0x00A8
    x"80",x"90",x"90",x"90",x"90",x"FD",x"FD",x"00", -- 0x00B0
    x"9D",x"9D",x"91",x"81",x"C5",x"7C",x"38",x"00", -- 0x00B8
    x"FD",x"FD",x"10",x"10",x"10",x"FD",x"FD",x"00", -- 0x00C0
    x"81",x"81",x"FD",x"FD",x"81",x"81",x"00",x"00", -- 0x00C8
    x"FC",x"FD",x"01",x"01",x"01",x"05",x"04",x"00", -- 0x00D0
    x"81",x"C5",x"6D",x"3C",x"18",x"FD",x"FD",x"00", -- 0x00D8
    x"01",x"01",x"01",x"01",x"FD",x"FD",x"00",x"00", -- 0x00E0
    x"FD",x"FD",x"70",x"38",x"70",x"FD",x"FD",x"00", -- 0x00E8
    x"FD",x"FD",x"1C",x"38",x"70",x"FD",x"FD",x"00", -- 0x00F0
    x"7C",x"FD",x"81",x"81",x"81",x"FD",x"7C",x"00", -- 0x00F8
    x"70",x"F8",x"88",x"88",x"88",x"FD",x"FD",x"00", -- 0x0100
    x"79",x"FC",x"8D",x"89",x"81",x"FD",x"7C",x"00", -- 0x0108
    x"71",x"F5",x"9D",x"8C",x"88",x"FD",x"FD",x"00", -- 0x0110
    x"0C",x"5D",x"D1",x"91",x"91",x"F5",x"64",x"00", -- 0x0118
    x"80",x"80",x"FD",x"FD",x"80",x"80",x"00",x"00", -- 0x0120
    x"FC",x"FD",x"01",x"01",x"01",x"FD",x"FC",x"00", -- 0x0128
    x"F0",x"F8",x"1C",x"0D",x"1C",x"F8",x"F0",x"00", -- 0x0130
    x"F8",x"FD",x"1C",x"38",x"1C",x"FD",x"F8",x"00", -- 0x0138
    x"C5",x"ED",x"7C",x"38",x"7C",x"ED",x"C5",x"00", -- 0x0140
    x"C0",x"F0",x"1D",x"1D",x"F0",x"C0",x"00",x"00", -- 0x0148
    x"C1",x"E1",x"F1",x"B9",x"9D",x"8D",x"85",x"00", -- 0x0150
    x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00", -- 0x0158
    x"00",x"00",x"00",x"00",x"08",x"0C",x"0D",x"0F", -- 0x0160
    x"00",x"00",x"80",x"00",x"08",x"18",x"38",x"78", -- 0x0168
    x"07",x"02",x"02",x"00",x"00",x"00",x"00",x"00", -- 0x0170
    x"70",x"40",x"C0",x"80",x"80",x"00",x"00",x"00", -- 0x0178
    x"04",x"0F",x"0F",x"0F",x"0F",x"0F",x"07",x"07", -- 0x0180
    x"20",x"F0",x"F0",x"F0",x"F0",x"F0",x"E0",x"E0", -- 0x0188
    x"0F",x"0F",x"0F",x"0F",x"0F",x"0E",x"07",x"00", -- 0x0190
    x"F0",x"F0",x"F0",x"F0",x"F0",x"B0",x"E0",x"00", -- 0x0198
    x"00",x"00",x"00",x"00",x"04",x"0C",x"00",x"00", -- 0x01A0
    x"00",x"00",x"80",x"00",x"10",x"58",x"20",x"10", -- 0x01A8
    x"00",x"00",x"00",x"0C",x"04",x"02",x"00",x"00", -- 0x01B0
    x"10",x"10",x"20",x"18",x"10",x"C0",x"80",x"00", -- 0x01B8
    x"00",x"02",x"00",x"08",x"18",x"0C",x"00",x"00", -- 0x01C0
    x"00",x"00",x"80",x"08",x"0C",x"58",x"20",x"10", -- 0x01C8
    x"00",x"00",x"00",x"0C",x"18",x"0A",x"02",x"00", -- 0x01D0
    x"10",x"10",x"20",x"18",x"0C",x"C8",x"C0",x"80", -- 0x01D8
    x"00",x"00",x"00",x"08",x"18",x"0C",x"00",x"00", -- 0x01E0
    x"00",x"40",x"80",x"08",x"0C",x"58",x"20",x"10", -- 0x01E8
    x"00",x"08",x"18",x"0C",x"00",x"02",x"02",x"00", -- 0x01F0
    x"10",x"18",x"2C",x"18",x"00",x"C0",x"C0",x"80", -- 0x01F8
    x"7E",x"D7",x"B3",x"F7",x"5F",x"CC",x"D8",x"F8", -- 0x0200
    x"FB",x"DA",x"9B",x"BF",x"FF",x"41",x"00",x"00", -- 0x0208
    x"E8",x"B8",x"98",x"BC",x"F8",x"10",x"00",x"00", -- 0x0210
    x"B8",x"9C",x"B8",x"F8",x"58",x"C8",x"DC",x"F8", -- 0x0218
    x"78",x"F8",x"DC",x"97",x"B3",x"F7",x"DF",x"76", -- 0x0220
    x"00",x"00",x"41",x"FF",x"F7",x"B3",x"97",x"BD", -- 0x0228
    x"00",x"00",x"10",x"F8",x"BD",x"98",x"B8",x"E8", -- 0x0230
    x"77",x"FE",x"BC",x"FE",x"EF",x"E7",x"EE",x"7F", -- 0x0238
    x"00",x"10",x"38",x"10",x"01",x"07",x"01",x"17", -- 0x0240
    x"00",x"00",x"20",x"70",x"20",x"00",x"08",x"AC", -- 0x0248
    x"3A",x"10",x"00",x"02",x"13",x"3A",x"10",x"00", -- 0x0250
    x"C8",x"80",x"04",x"0D",x"84",x"12",x"38",x"10", -- 0x0258
    x"00",x"1C",x"3D",x"1D",x"3D",x"1C",x"00",x"00", -- 0x0260
    x"67",x"3C",x"3C",x"7C",x"3C",x"3C",x"67",x"00", -- 0x0268
    x"3C",x"41",x"82",x"A6",x"A6",x"9A",x"41",x"3C", -- 0x0270
    x"FF",x"82",x"82",x"82",x"82",x"82",x"82",x"FF", -- 0x0278
    x"01",x"03",x"05",x"0F",x"05",x"07",x"05",x"07", -- 0x0280
    x"40",x"C0",x"60",x"F0",x"60",x"E0",x"60",x"E0", -- 0x0288
    x"07",x"07",x"07",x"0F",x"07",x"07",x"03",x"02", -- 0x0290
    x"E0",x"E0",x"E0",x"F0",x"E0",x"E0",x"C0",x"80", -- 0x0298
    x"02",x"02",x"00",x"00",x"00",x"08",x"00",x"00", -- 0x02A0
    x"38",x"38",x"38",x"38",x"D0",x"18",x"18",x"18", -- 0x02A8
    x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B0
    x"00",x"90",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"01",x"00",x"00",x"00",x"04",x"04",x"00", -- 0x02C0
    x"38",x"18",x"18",x"58",x"50",x"58",x"18",x"38", -- 0x02C8
    x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"08", -- 0x02D0
    x"38",x"38",x"38",x"38",x"30",x"B8",x"38",x"38", -- 0x02D8
    x"00",x"00",x"00",x"03",x"0D",x"18",x"18",x"18", -- 0x02E0
    x"00",x"00",x"00",x"C0",x"70",x"18",x"C8",x"00", -- 0x02E8
    x"0D",x"02",x"00",x"08",x"00",x"00",x"00",x"00", -- 0x02F0
    x"78",x"F8",x"78",x"30",x"78",x"78",x"38",x"38", -- 0x02F8
    x"07",x"08",x"08",x"08",x"07",x"00",x"07",x"08", -- 0x0300
    x"C0",x"20",x"20",x"20",x"C0",x"00",x"C0",x"20", -- 0x0308
    x"08",x"08",x"07",x"00",x"00",x"0F",x"04",x"00", -- 0x0310
    x"20",x"20",x"C0",x"00",x"20",x"E0",x"20",x"00", -- 0x0318
    x"07",x"08",x"08",x"07",x"00",x"07",x"08",x"08", -- 0x0320
    x"C0",x"20",x"20",x"C0",x"00",x"C0",x"20",x"20", -- 0x0328
    x"07",x"00",x"05",x"0A",x"08",x"08",x"04",x"00", -- 0x0330
    x"C0",x"00",x"20",x"20",x"A0",x"60",x"20",x"00", -- 0x0338
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0340
    x"00",x"20",x"20",x"20",x"20",x"21",x"26",x"22", -- 0x0348
    x"00",x"00",x"00",x"00",x"03",x"03",x"00",x"00", -- 0x0350
    x"40",x"41",x"06",x"02",x"02",x"02",x"42",x"20", -- 0x0358
    x"02",x"03",x"62",x"90",x"97",x"7F",x"3B",x"3E", -- 0x0360
    x"E0",x"FA",x"FB",x"FF",x"FD",x"FF",x"FC",x"E4", -- 0x0368
    x"3E",x"3B",x"7F",x"97",x"90",x"62",x"03",x"02", -- 0x0370
    x"E4",x"E4",x"FF",x"FD",x"FF",x"FB",x"FA",x"E0", -- 0x0378
    x"00",x"00",x"10",x"3C",x"01",x"07",x"1F",x"1F", -- 0x0380
    x"00",x"00",x"04",x"1D",x"30",x"E0",x"E0",x"E0", -- 0x0388
    x"1F",x"1F",x"07",x"01",x"3C",x"10",x"00",x"00", -- 0x0390
    x"E0",x"E0",x"E0",x"30",x"1D",x"04",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"10",x"3D",x"07",x"1F",x"1F", -- 0x03A0
    x"00",x"00",x"00",x"10",x"38",x"EC",x"E3",x"E0", -- 0x03A8
    x"1F",x"1F",x"07",x"3D",x"10",x"00",x"00",x"00", -- 0x03B0
    x"E0",x"E3",x"EC",x"38",x"10",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"08",x"1D",x"01",x"07",x"1F",x"1F", -- 0x03C0
    x"00",x"00",x"20",x"F0",x"80",x"C0",x"E0",x"E0", -- 0x03C8
    x"1F",x"1F",x"07",x"01",x"1D",x"08",x"00",x"00", -- 0x03D0
    x"E0",x"E0",x"C0",x"80",x"F0",x"20",x"00",x"00", -- 0x03D8
    x"00",x"10",x"30",x"10",x"18",x"0F",x"07",x"07", -- 0x03E0
    x"00",x"08",x"0C",x"08",x"18",x"F0",x"E0",x"E0", -- 0x03E8
    x"07",x"0F",x"17",x"13",x"33",x"10",x"00",x"00", -- 0x03F0
    x"E0",x"F0",x"E8",x"C8",x"CC",x"08",x"00",x"00", -- 0x03F8
    x"00",x"01",x"05",x"0C",x"18",x"0F",x"07",x"07", -- 0x0400
    x"00",x"40",x"60",x"30",x"18",x"F0",x"E0",x"E0", -- 0x0408
    x"07",x"0F",x"0F",x"0B",x"1B",x"08",x"00",x"00", -- 0x0410
    x"E0",x"F0",x"F0",x"D0",x"D8",x"10",x"00",x"00", -- 0x0418
    x"00",x"00",x"00",x"00",x"10",x"33",x"17",x"1F", -- 0x0420
    x"00",x"00",x"00",x"00",x"08",x"CC",x"E8",x"F8", -- 0x0428
    x"07",x"1F",x"17",x"33",x"13",x"00",x"00",x"00", -- 0x0430
    x"E0",x"F8",x"E8",x"CC",x"C8",x"00",x"00",x"00", -- 0x0438
    x"00",x"00",x"01",x"08",x"12",x"07",x"27",x"0F", -- 0x0440
    x"00",x"00",x"40",x"10",x"88",x"E0",x"E4",x"F0", -- 0x0448
    x"0F",x"27",x"07",x"12",x"08",x"01",x"00",x"00", -- 0x0450
    x"F0",x"E4",x"E0",x"88",x"10",x"40",x"00",x"00", -- 0x0458
    x"00",x"02",x"14",x"20",x"02",x"46",x"03",x"4F", -- 0x0460
    x"00",x"80",x"28",x"04",x"80",x"A1",x"C0",x"F1", -- 0x0468
    x"4F",x"03",x"46",x"02",x"20",x"14",x"02",x"00", -- 0x0470
    x"F1",x"C0",x"A1",x"80",x"04",x"28",x"80",x"00", -- 0x0478
    x"01",x"00",x"20",x"00",x"01",x"00",x"88",x"02", -- 0x0480
    x"40",x"00",x"04",x"00",x"40",x"00",x"12",x"80", -- 0x0488
    x"02",x"88",x"00",x"01",x"00",x"20",x"00",x"01", -- 0x0490
    x"80",x"12",x"00",x"40",x"00",x"04",x"00",x"40", -- 0x0498
    x"00",x"00",x"00",x"04",x"0A",x"03",x"07",x"07", -- 0x04A0
    x"00",x"00",x"00",x"10",x"88",x"C0",x"E0",x"E0", -- 0x04A8
    x"07",x"07",x"03",x"12",x"08",x"00",x"00",x"00", -- 0x04B0
    x"E0",x"E0",x"C0",x"88",x"10",x"00",x"00",x"00", -- 0x04B8
    x"00",x"02",x"00",x"00",x"00",x"01",x"04",x"22", -- 0x04C0
    x"00",x"80",x"00",x"00",x"00",x"20",x"90",x"C1", -- 0x04C8
    x"22",x"02",x"04",x"01",x"00",x"00",x"02",x"00", -- 0x04D0
    x"C1",x"C0",x"90",x"20",x"00",x"00",x"80",x"00", -- 0x04D8
    x"02",x"00",x"00",x"01",x"01",x"00",x"00",x"00", -- 0x04E0
    x"00",x"08",x"14",x"01",x"21",x"29",x"48",x"48", -- 0x04E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F0
    x"08",x"00",x"04",x"04",x"06",x"02",x"0A",x"08", -- 0x04F8
    x"02",x"03",x"07",x"07",x"0F",x"07",x"07",x"07", -- 0x0500
    x"80",x"C0",x"E0",x"E0",x"F0",x"E0",x"E0",x"E0", -- 0x0508
    x"07",x"05",x"05",x"05",x"0F",x"05",x"05",x"01", -- 0x0510
    x"E0",x"60",x"E0",x"60",x"F0",x"60",x"E0",x"40", -- 0x0518
    x"00",x"29",x"29",x"3F",x"08",x"08",x"0F",x"07", -- 0x0520
    x"00",x"54",x"54",x"FC",x"10",x"10",x"F0",x"E0", -- 0x0528
    x"07",x"3F",x"07",x"37",x"07",x"3F",x"03",x"00", -- 0x0530
    x"EC",x"F0",x"EC",x"E0",x"EC",x"F0",x"CC",x"00", -- 0x0538
    x"0F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"1F", -- 0x0540
    x"F0",x"F0",x"F8",x"F8",x"F8",x"F0",x"00",x"F8", -- 0x0548
    x"1F",x"1F",x"0F",x"07",x"00",x"00",x"00",x"00", -- 0x0550
    x"F8",x"F8",x"F0",x"E0",x"00",x"00",x"00",x"00", -- 0x0558
    x"00",x"00",x"0F",x"1F",x"1F",x"1F",x"0F",x"0F", -- 0x0560
    x"00",x"00",x"F0",x"F8",x"F8",x"F8",x"F0",x"F0", -- 0x0568
    x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x0570
    x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x0578
    x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00", -- 0x0580
    x"20",x"08",x"00",x"10",x"00",x"40",x"00",x"00", -- 0x0588
    x"00",x"00",x"21",x"02",x"00",x"00",x"00",x"00", -- 0x0590
    x"00",x"00",x"00",x"00",x"80",x"40",x"00",x"00", -- 0x0598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A0
    x"00",x"10",x"00",x"00",x"08",x"00",x"00",x"10", -- 0x05A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B0
    x"00",x"40",x"00",x"00",x"40",x"00",x"10",x"00", -- 0x05B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C0
    x"00",x"20",x"00",x"00",x"10",x"00",x"20",x"00", -- 0x05C8
    x"00",x"00",x"00",x"08",x"00",x"00",x"00",x"00", -- 0x05D0
    x"80",x"00",x"00",x"80",x"80",x"80",x"00",x"00", -- 0x05D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E0
    x"00",x"00",x"20",x"00",x"00",x"00",x"40",x"00", -- 0x05E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F0
    x"80",x"00",x"00",x"40",x"00",x"00",x"20",x"08", -- 0x05F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0600
    x"80",x"00",x"20",x"00",x"00",x"10",x"00",x"08", -- 0x0608
    x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00", -- 0x0610
    x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0618
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0620
    x"00",x"00",x"00",x"80",x"00",x"00",x"40",x"00", -- 0x0628
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0630
    x"00",x"08",x"00",x"00",x"10",x"00",x"20",x"00", -- 0x0638
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0640
    x"02",x"02",x"66",x"06",x"04",x"44",x"10",x"00", -- 0x0648
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0650
    x"21",x"81",x"09",x"49",x"09",x"08",x"10",x"10", -- 0x0658
    x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x0660
    x"02",x"02",x"84",x"04",x"00",x"21",x"46",x"02", -- 0x0668
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0670
    x"86",x"02",x"0A",x"0A",x"40",x"44",x"14",x"14", -- 0x0678
    x"00",x"00",x"00",x"00",x"18",x"00",x"0C",x"00", -- 0x0680
    x"00",x"00",x"20",x"00",x"20",x"01",x"46",x"02", -- 0x0688
    x"03",x"00",x"00",x"00",x"05",x"05",x"00",x"00", -- 0x0690
    x"60",x"01",x"06",x"02",x"02",x"C2",x"82",x"20", -- 0x0698
    x"C0",x"E0",x"E3",x"E3",x"E3",x"E3",x"E3",x"E3", -- 0x06A0
    x"00",x"00",x"00",x"80",x"80",x"80",x"80",x"80", -- 0x06A8
    x"E3",x"E3",x"FF",x"FF",x"FF",x"FF",x"00",x"00", -- 0x06B0
    x"80",x"80",x"FC",x"FD",x"FD",x"FD",x"01",x"00", -- 0x06B8
    x"7F",x"7F",x"FF",x"FF",x"C3",x"E3",x"E0",x"E0", -- 0x06C0
    x"0C",x"8D",x"BD",x"BD",x"FD",x"FD",x"F1",x"F8", -- 0x06C8
    x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"00",x"00", -- 0x06D0
    x"F8",x"F8",x"FC",x"FD",x"FD",x"FD",x"01",x"00", -- 0x06D8
    x"3F",x"3F",x"FF",x"FF",x"C0",x"E0",x"E0",x"E0", -- 0x06E0
    x"F0",x"F8",x"FC",x"FD",x"0D",x"0D",x"0D",x"0D", -- 0x06E8
    x"E0",x"E0",x"FF",x"FF",x"3F",x"3F",x"00",x"00", -- 0x06F0
    x"0D",x"0D",x"FD",x"FD",x"F1",x"F8",x"08",x"00", -- 0x06F8
    x"00",x"00",x"08",x"40",x"48",x"00",x"00",x"00", -- 0x0700
    x"00",x"08",x"04",x"31",x"29",x"49",x"28",x"0A", -- 0x0708
    x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"02", -- 0x0710
    x"2A",x"02",x"16",x"14",x"14",x"14",x"04",x"20", -- 0x0718
    x"00",x"00",x"10",x"3B",x"7F",x"33",x"13",x"1F", -- 0x0720
    x"00",x"00",x"08",x"DC",x"FD",x"FC",x"F8",x"F8", -- 0x0728
    x"1F",x"13",x"33",x"7F",x"3B",x"10",x"00",x"00", -- 0x0730
    x"F8",x"FC",x"FD",x"DC",x"08",x"00",x"00",x"00", -- 0x0738
    x"00",x"30",x"77",x"7F",x"33",x"37",x"7F",x"7F", -- 0x0740
    x"00",x"18",x"D8",x"FC",x"FC",x"F8",x"F8",x"F8", -- 0x0748
    x"7F",x"7F",x"37",x"33",x"7F",x"77",x"30",x"00", -- 0x0750
    x"F8",x"F8",x"F8",x"FC",x"FC",x"D8",x"18",x"00", -- 0x0758
    x"30",x"63",x"FF",x"F8",x"BC",x"7F",x"7F",x"7F", -- 0x0760
    x"0C",x"CC",x"FF",x"FF",x"FE",x"FD",x"FD",x"FD", -- 0x0768
    x"7F",x"7F",x"7F",x"BC",x"F8",x"FF",x"63",x"30", -- 0x0770
    x"FD",x"FD",x"FD",x"FE",x"FF",x"FF",x"CC",x"00", -- 0x0778
    x"0C",x"0C",x"01",x"3A",x"68",x"DC",x"FD",x"FD", -- 0x0780
    x"00",x"00",x"00",x"03",x"83",x"44",x"28",x"10", -- 0x0788
    x"FD",x"DC",x"68",x"3A",x"01",x"0C",x"0C",x"00", -- 0x0790
    x"28",x"44",x"83",x"03",x"00",x"00",x"00",x"00", -- 0x0798
    x"C3",x"E3",x"E3",x"E3",x"E3",x"E3",x"E0",x"E0", -- 0x07A0
    x"FC",x"FD",x"FD",x"FD",x"0D",x"8D",x"8D",x"0D", -- 0x07A8
    x"F0",x"F8",x"3F",x"3F",x"0F",x"0F",x"00",x"00", -- 0x07B0
    x"3D",x"3D",x"F1",x"F8",x"C8",x"E0",x"20",x"00", -- 0x07B8
    x"C0",x"E0",x"E3",x"E3",x"E3",x"E3",x"E3",x"E3", -- 0x07C0
    x"0C",x"0D",x"0D",x"8D",x"8D",x"8D",x"8D",x"8D", -- 0x07C8
    x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x07D0
    x"FD",x"FD",x"FD",x"FD",x"01",x"00",x"00",x"00", -- 0x07D8
    x"02",x"03",x"62",x"90",x"97",x"7F",x"3A",x"38", -- 0x07E0
    x"E0",x"FA",x"FB",x"FF",x"FD",x"FF",x"FC",x"E4", -- 0x07E8
    x"38",x"3A",x"7F",x"97",x"90",x"62",x"03",x"02", -- 0x07F0
    x"E4",x"E4",x"FF",x"FD",x"FF",x"FB",x"FA",x"E0"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
