library work;
use work.pace_pkg.all;
use work.project_pkg.all;

package body platform_pkg is

    constant CABAL_SRC_DIR    : string := "../../../../../src/platform/cabal/";

end platform_pkg;
