-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_SND_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_SND_1 is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"0C",x"80",x"77",x"C9",x"B7",x"C8",x"21",x"17", -- 0x0000
    x"08",x"E5",x"87",x"5F",x"16",x"00",x"21",x"60", -- 0x0008
    x"08",x"19",x"5E",x"23",x"56",x"EB",x"E9",x"B7", -- 0x0010
    x"C8",x"3A",x"10",x"80",x"FE",x"01",x"28",x"18", -- 0x0018
    x"FE",x"02",x"28",x"1C",x"FE",x"03",x"28",x"20", -- 0x0020
    x"FE",x"04",x"28",x"24",x"FE",x"05",x"28",x"28", -- 0x0028
    x"AF",x"32",x"0A",x"80",x"32",x"0B",x"80",x"C9", -- 0x0030
    x"AF",x"32",x"00",x"80",x"32",x"01",x"80",x"C9", -- 0x0038
    x"AF",x"32",x"02",x"80",x"32",x"03",x"80",x"C9", -- 0x0040
    x"AF",x"32",x"04",x"80",x"32",x"05",x"80",x"C9", -- 0x0048
    x"AF",x"32",x"06",x"80",x"32",x"07",x"80",x"C9", -- 0x0050
    x"AF",x"32",x"08",x"80",x"32",x"09",x"80",x"C9", -- 0x0058
    x"00",x"00",x"39",x"09",x"B5",x"09",x"31",x"0A", -- 0x0060
    x"AD",x"0A",x"29",x"0B",x"1F",x"0D",x"4E",x"12", -- 0x0068
    x"CE",x"13",x"CE",x"0D",x"D4",x"0D",x"4A",x"10", -- 0x0070
    x"51",x"10",x"58",x"10",x"C7",x"10",x"CE",x"10", -- 0x0078
    x"00",x"00",x"00",x"00",x"20",x"11",x"73",x"0B", -- 0x0080
    x"12",x"0C",x"A3",x"0C",x"00",x"00",x"00",x"00", -- 0x0088
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0098
    x"97",x"0D",x"B1",x"11",x"1A",x"12",x"DE",x"12", -- 0x00A0
    x"5B",x"13",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B8
    x"CD",x"2C",x"0B",x"3E",x"03",x"32",x"1B",x"80", -- 0x00C0
    x"3E",x"0F",x"32",x"1C",x"80",x"3E",x"1F",x"32", -- 0x00C8
    x"1D",x"80",x"21",x"80",x"00",x"22",x"1E",x"80", -- 0x00D0
    x"22",x"20",x"80",x"3E",x"04",x"32",x"22",x"80", -- 0x00D8
    x"3E",x"40",x"32",x"23",x"80",x"32",x"24",x"80", -- 0x00E0
    x"3E",x"03",x"32",x"26",x"80",x"3E",x"0A",x"32", -- 0x00E8
    x"27",x"80",x"21",x"00",x"08",x"22",x"28",x"80", -- 0x00F0
    x"3E",x"08",x"32",x"2A",x"80",x"32",x"2B",x"80", -- 0x00F8
    x"21",x"40",x"00",x"22",x"2C",x"80",x"22",x"2E", -- 0x0100
    x"80",x"3E",x"0C",x"32",x"30",x"80",x"3E",x"03", -- 0x0108
    x"32",x"32",x"80",x"3E",x"0A",x"32",x"33",x"80", -- 0x0110
    x"21",x"00",x"02",x"22",x"34",x"80",x"21",x"00", -- 0x0118
    x"08",x"22",x"36",x"80",x"21",x"00",x"02",x"22", -- 0x0120
    x"38",x"80",x"3E",x"08",x"32",x"3A",x"80",x"32", -- 0x0128
    x"3B",x"80",x"21",x"20",x"00",x"22",x"3D",x"80", -- 0x0130
    x"C9",x"3E",x"FF",x"C9",x"CD",x"2C",x"0B",x"3E", -- 0x0138
    x"03",x"32",x"1B",x"80",x"3E",x"0F",x"32",x"1C", -- 0x0140
    x"80",x"3E",x"1F",x"32",x"1D",x"80",x"21",x"80", -- 0x0148
    x"00",x"22",x"1E",x"80",x"22",x"20",x"80",x"3E", -- 0x0150
    x"01",x"32",x"22",x"80",x"3E",x"20",x"32",x"23", -- 0x0158
    x"80",x"32",x"24",x"80",x"3E",x"03",x"32",x"26", -- 0x0160
    x"80",x"3E",x"0D",x"32",x"27",x"80",x"21",x"00", -- 0x0168
    x"08",x"22",x"28",x"80",x"3E",x"08",x"32",x"2A", -- 0x0170
    x"80",x"32",x"2B",x"80",x"21",x"40",x"00",x"22", -- 0x0178
    x"2C",x"80",x"22",x"2E",x"80",x"3E",x"02",x"32", -- 0x0180
    x"30",x"80",x"3E",x"03",x"32",x"32",x"80",x"3E", -- 0x0188
    x"0E",x"32",x"33",x"80",x"21",x"00",x"02",x"22", -- 0x0190
    x"34",x"80",x"21",x"00",x"08",x"22",x"36",x"80", -- 0x0198
    x"21",x"01",x"00",x"22",x"38",x"80",x"3E",x"18", -- 0x01A0
    x"32",x"3A",x"80",x"32",x"3B",x"80",x"21",x"00", -- 0x01A8
    x"01",x"22",x"3D",x"80",x"C9",x"3E",x"FF",x"C9", -- 0x01B0
    x"CD",x"2C",x"0B",x"3E",x"02",x"32",x"1B",x"80", -- 0x01B8
    x"3E",x"0F",x"32",x"1C",x"80",x"3E",x"08",x"32", -- 0x01C0
    x"1D",x"80",x"21",x"80",x"00",x"22",x"1E",x"80", -- 0x01C8
    x"22",x"20",x"80",x"3E",x"01",x"32",x"22",x"80", -- 0x01D0
    x"3E",x"20",x"32",x"23",x"80",x"32",x"24",x"80", -- 0x01D8
    x"3E",x"03",x"32",x"26",x"80",x"3E",x"0A",x"32", -- 0x01E0
    x"27",x"80",x"21",x"00",x"08",x"22",x"28",x"80", -- 0x01E8
    x"3E",x"08",x"32",x"2A",x"80",x"32",x"2B",x"80", -- 0x01F0
    x"21",x"40",x"00",x"22",x"2C",x"80",x"22",x"2E", -- 0x01F8
    x"80",x"3E",x"03",x"32",x"30",x"80",x"3E",x"03", -- 0x0200
    x"32",x"32",x"80",x"3E",x"08",x"32",x"33",x"80", -- 0x0208
    x"21",x"00",x"02",x"22",x"34",x"80",x"21",x"00", -- 0x0210
    x"08",x"22",x"36",x"80",x"21",x"01",x"00",x"22", -- 0x0218
    x"38",x"80",x"3E",x"20",x"32",x"3A",x"80",x"32", -- 0x0220
    x"3B",x"80",x"21",x"20",x"00",x"22",x"3D",x"80", -- 0x0228
    x"C9",x"3E",x"FF",x"C9",x"CD",x"2C",x"0B",x"3E", -- 0x0230
    x"03",x"32",x"1B",x"80",x"3E",x"0E",x"32",x"1C", -- 0x0238
    x"80",x"3E",x"1F",x"32",x"1D",x"80",x"21",x"80", -- 0x0240
    x"00",x"22",x"1E",x"80",x"22",x"20",x"80",x"3E", -- 0x0248
    x"01",x"32",x"22",x"80",x"3E",x"20",x"32",x"23", -- 0x0250
    x"80",x"32",x"24",x"80",x"3E",x"03",x"32",x"26", -- 0x0258
    x"80",x"3E",x"0C",x"32",x"27",x"80",x"21",x"00", -- 0x0260
    x"08",x"22",x"28",x"80",x"3E",x"08",x"32",x"2A", -- 0x0268
    x"80",x"32",x"2B",x"80",x"21",x"40",x"00",x"22", -- 0x0270
    x"2C",x"80",x"22",x"2E",x"80",x"3E",x"03",x"32", -- 0x0278
    x"30",x"80",x"3E",x"03",x"32",x"32",x"80",x"3E", -- 0x0280
    x"0F",x"32",x"33",x"80",x"21",x"00",x"02",x"22", -- 0x0288
    x"34",x"80",x"21",x"00",x"08",x"22",x"36",x"80", -- 0x0290
    x"21",x"01",x"00",x"22",x"38",x"80",x"3E",x"20", -- 0x0298
    x"32",x"3A",x"80",x"32",x"3B",x"80",x"21",x"20", -- 0x02A0
    x"00",x"22",x"3D",x"80",x"C9",x"3E",x"FF",x"C9", -- 0x02A8
    x"CD",x"2C",x"0B",x"3E",x"03",x"32",x"1B",x"80", -- 0x02B0
    x"3E",x"0F",x"32",x"1C",x"80",x"3E",x"1F",x"32", -- 0x02B8
    x"1D",x"80",x"21",x"80",x"00",x"22",x"1E",x"80", -- 0x02C0
    x"22",x"20",x"80",x"3E",x"04",x"32",x"22",x"80", -- 0x02C8
    x"3E",x"40",x"32",x"23",x"80",x"32",x"24",x"80", -- 0x02D0
    x"3E",x"03",x"32",x"26",x"80",x"3E",x"0C",x"32", -- 0x02D8
    x"27",x"80",x"21",x"00",x"08",x"22",x"28",x"80", -- 0x02E0
    x"3E",x"08",x"32",x"2A",x"80",x"32",x"2B",x"80", -- 0x02E8
    x"21",x"30",x"00",x"22",x"2C",x"80",x"22",x"2E", -- 0x02F0
    x"80",x"3E",x"08",x"32",x"30",x"80",x"3E",x"03", -- 0x02F8
    x"32",x"32",x"80",x"3E",x"09",x"32",x"33",x"80", -- 0x0300
    x"21",x"00",x"02",x"22",x"34",x"80",x"21",x"00", -- 0x0308
    x"08",x"22",x"36",x"80",x"21",x"00",x"01",x"22", -- 0x0310
    x"38",x"80",x"3E",x"01",x"32",x"3A",x"80",x"32", -- 0x0318
    x"3B",x"80",x"21",x"20",x"00",x"22",x"3D",x"80", -- 0x0320
    x"C9",x"3E",x"FF",x"C9",x"3E",x"13",x"CD",x"6F", -- 0x0328
    x"00",x"3E",x"14",x"CD",x"6F",x"00",x"3E",x"15", -- 0x0330
    x"CD",x"6F",x"00",x"C9",x"3A",x"1B",x"80",x"FE", -- 0x0338
    x"00",x"28",x"21",x"FE",x"01",x"28",x"22",x"FE", -- 0x0340
    x"02",x"28",x"23",x"CD",x"BC",x"07",x"AF",x"32", -- 0x0348
    x"25",x"80",x"16",x"06",x"21",x"1D",x"80",x"5E", -- 0x0350
    x"CD",x"4C",x"05",x"CD",x"80",x"05",x"06",x"00", -- 0x0358
    x"CD",x"FE",x"05",x"C9",x"CD",x"C7",x"06",x"18", -- 0x0360
    x"E5",x"CD",x"48",x"07",x"18",x"E0",x"CD",x"82", -- 0x0368
    x"07",x"18",x"DB",x"16",x"06",x"21",x"1D",x"80", -- 0x0370
    x"5E",x"CD",x"4C",x"05",x"3A",x"25",x"80",x"FE", -- 0x0378
    x"00",x"28",x"1E",x"FE",x"01",x"28",x"27",x"FE", -- 0x0380
    x"02",x"28",x"3C",x"21",x"24",x"80",x"35",x"20", -- 0x0388
    x"0E",x"3A",x"23",x"80",x"77",x"CD",x"4B",x"06", -- 0x0390
    x"3D",x"28",x"3E",x"47",x"CD",x"FE",x"05",x"AF", -- 0x0398
    x"C9",x"3A",x"1C",x"80",x"47",x"CD",x"FE",x"05", -- 0x03A0
    x"21",x"25",x"80",x"34",x"18",x"DD",x"2A",x"20", -- 0x03A8
    x"80",x"2B",x"7C",x"B5",x"20",x"0C",x"2A",x"1E", -- 0x03B0
    x"80",x"22",x"20",x"80",x"21",x"25",x"80",x"34", -- 0x03B8
    x"18",x"C9",x"22",x"20",x"80",x"18",x"C4",x"21", -- 0x03C0
    x"22",x"80",x"35",x"20",x"06",x"21",x"25",x"80", -- 0x03C8
    x"34",x"18",x"B8",x"AF",x"32",x"25",x"80",x"18", -- 0x03D0
    x"B2",x"16",x"06",x"1E",x"04",x"CD",x"4C",x"05", -- 0x03D8
    x"3E",x"FF",x"C9",x"3A",x"26",x"80",x"FE",x"00", -- 0x03E0
    x"28",x"19",x"FE",x"01",x"28",x"1A",x"FE",x"02", -- 0x03E8
    x"28",x"1B",x"CD",x"BC",x"07",x"AF",x"32",x"31", -- 0x03F0
    x"80",x"2A",x"28",x"80",x"CD",x"C6",x"04",x"CD", -- 0x03F8
    x"0D",x"05",x"C9",x"CD",x"C7",x"06",x"18",x"ED", -- 0x0400
    x"CD",x"48",x"07",x"18",x"E8",x"CD",x"82",x"07", -- 0x0408
    x"18",x"E3",x"3A",x"31",x"80",x"FE",x"00",x"28", -- 0x0410
    x"1F",x"FE",x"01",x"28",x"2E",x"2A",x"2E",x"80", -- 0x0418
    x"2B",x"7C",x"B5",x"20",x"40",x"2A",x"2C",x"80", -- 0x0420
    x"22",x"2E",x"80",x"21",x"30",x"80",x"35",x"28", -- 0x0428
    x"39",x"21",x"31",x"80",x"36",x"00",x"AF",x"C9", -- 0x0430
    x"3A",x"27",x"80",x"47",x"CD",x"FE",x"05",x"3A", -- 0x0438
    x"2A",x"80",x"32",x"2B",x"80",x"21",x"31",x"80", -- 0x0440
    x"34",x"18",x"EB",x"21",x"2B",x"80",x"35",x"20", -- 0x0448
    x"CC",x"3A",x"2A",x"80",x"77",x"CD",x"4B",x"06", -- 0x0450
    x"3D",x"20",x"04",x"21",x"31",x"80",x"34",x"47", -- 0x0458
    x"CD",x"FE",x"05",x"18",x"B8",x"22",x"2E",x"80", -- 0x0460
    x"18",x"CC",x"3E",x"FF",x"C9",x"3A",x"32",x"80", -- 0x0468
    x"FE",x"00",x"28",x"20",x"FE",x"01",x"28",x"21", -- 0x0470
    x"FE",x"02",x"28",x"22",x"CD",x"BC",x"07",x"AF", -- 0x0478
    x"32",x"3C",x"80",x"2A",x"36",x"80",x"CD",x"C6", -- 0x0480
    x"04",x"CD",x"0D",x"05",x"3A",x"33",x"80",x"47", -- 0x0488
    x"CD",x"FE",x"05",x"C9",x"CD",x"C7",x"06",x"18", -- 0x0490
    x"E6",x"CD",x"48",x"07",x"18",x"E1",x"CD",x"82", -- 0x0498
    x"07",x"18",x"DC",x"3A",x"3C",x"80",x"FE",x"00", -- 0x04A0
    x"28",x"22",x"FE",x"01",x"28",x"32",x"CD",x"80", -- 0x04A8
    x"06",x"B7",x"ED",x"5B",x"3D",x"80",x"ED",x"52", -- 0x04B0
    x"ED",x"5B",x"34",x"80",x"7C",x"BA",x"20",x"07", -- 0x04B8
    x"7D",x"BB",x"20",x"03",x"2A",x"36",x"80",x"CD", -- 0x04C0
    x"C6",x"04",x"AF",x"C9",x"2A",x"38",x"80",x"2B", -- 0x04C8
    x"7C",x"B5",x"20",x"07",x"3E",x"01",x"32",x"3C", -- 0x04D0
    x"80",x"18",x"D3",x"22",x"38",x"80",x"18",x"CE", -- 0x04D8
    x"21",x"3A",x"80",x"35",x"20",x"C8",x"3A",x"3B", -- 0x04E0
    x"80",x"77",x"CD",x"4B",x"06",x"3D",x"28",x"06", -- 0x04E8
    x"47",x"CD",x"FE",x"05",x"18",x"B8",x"3E",x"FF", -- 0x04F0
    x"C9",x"CD",x"48",x"07",x"AF",x"32",x"43",x"80", -- 0x04F8
    x"3E",x"02",x"32",x"42",x"80",x"CD",x"0D",x"05", -- 0x0500
    x"3E",x"08",x"32",x"3F",x"80",x"21",x"20",x"00", -- 0x0508
    x"22",x"40",x"80",x"21",x"40",x"00",x"CD",x"C6", -- 0x0510
    x"04",x"06",x"08",x"CD",x"FE",x"05",x"C9",x"3A", -- 0x0518
    x"43",x"80",x"B7",x"20",x"0B",x"2A",x"40",x"80", -- 0x0520
    x"2B",x"7C",x"B5",x"28",x"37",x"22",x"40",x"80", -- 0x0528
    x"21",x"3F",x"80",x"35",x"28",x"1A",x"CD",x"80", -- 0x0530
    x"06",x"11",x"10",x"00",x"19",x"11",x"00",x"02", -- 0x0538
    x"7C",x"BA",x"20",x"07",x"7D",x"BB",x"20",x"03", -- 0x0540
    x"21",x"40",x"00",x"CD",x"C6",x"04",x"AF",x"C9", -- 0x0548
    x"3E",x"08",x"32",x"3F",x"80",x"CD",x"4B",x"06", -- 0x0550
    x"3D",x"28",x"06",x"47",x"CD",x"FE",x"05",x"18", -- 0x0558
    x"D5",x"3E",x"FF",x"C9",x"21",x"20",x"00",x"22", -- 0x0560
    x"40",x"80",x"21",x"42",x"80",x"35",x"20",x"05", -- 0x0568
    x"3E",x"01",x"32",x"43",x"80",x"CD",x"08",x"0D", -- 0x0570
    x"18",x"A5",x"CD",x"82",x"07",x"3E",x"08",x"32", -- 0x0578
    x"44",x"80",x"21",x"00",x"0A",x"22",x"45",x"80", -- 0x0580
    x"21",x"40",x"00",x"CD",x"C6",x"04",x"CD",x"0D", -- 0x0588
    x"05",x"06",x"0B",x"CD",x"FE",x"05",x"C9",x"2A", -- 0x0590
    x"45",x"80",x"2B",x"7C",x"B5",x"28",x"17",x"22", -- 0x0598
    x"45",x"80",x"21",x"44",x"80",x"35",x"20",x"0C", -- 0x05A0
    x"36",x"08",x"CD",x"80",x"06",x"11",x"02",x"00", -- 0x05A8
    x"19",x"CD",x"C6",x"04",x"AF",x"C9",x"3E",x"FF", -- 0x05B0
    x"C9",x"CD",x"C7",x"06",x"3E",x"00",x"32",x"73", -- 0x05B8
    x"80",x"CD",x"0D",x"05",x"C3",x"8E",x"0F",x"CD", -- 0x05C0
    x"C7",x"06",x"CD",x"0D",x"05",x"C9",x"DD",x"21", -- 0x05C8
    x"50",x"80",x"18",x"06",x"DD",x"21",x"58",x"80", -- 0x05D0
    x"18",x"00",x"DD",x"7E",x"00",x"FE",x"FF",x"C8", -- 0x05D8
    x"CD",x"E5",x"0D",x"AF",x"C9",x"DD",x"35",x"01", -- 0x05E0
    x"C0",x"3A",x"72",x"80",x"DD",x"77",x"01",x"DD", -- 0x05E8
    x"CB",x"00",x"46",x"C2",x"05",x"0E",x"DD",x"7E", -- 0x05F0
    x"07",x"D6",x"01",x"FA",x"05",x"0E",x"DD",x"77", -- 0x05F8
    x"07",x"47",x"CD",x"FE",x"05",x"DD",x"35",x"00", -- 0x0600
    x"C0",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"7E", -- 0x0608
    x"47",x"E6",x"1F",x"CA",x"9A",x"0E",x"FE",x"1F", -- 0x0610
    x"C2",x"B6",x"0E",x"23",x"DD",x"75",x"02",x"DD", -- 0x0618
    x"74",x"03",x"78",x"E6",x"E0",x"0F",x"0F",x"0F", -- 0x0620
    x"0F",x"4F",x"06",x"00",x"21",x"35",x"0E",x"09", -- 0x0628
    x"5E",x"23",x"56",x"D5",x"C9",x"45",x"0E",x"5D", -- 0x0630
    x"0E",x"73",x"0E",x"90",x"0E",x"90",x"0E",x"90", -- 0x0638
    x"0E",x"90",x"0E",x"90",x"0E",x"DD",x"6E",x"02", -- 0x0640
    x"DD",x"66",x"03",x"4E",x"CB",x"21",x"06",x"00", -- 0x0648
    x"21",x"E6",x"0E",x"09",x"5E",x"23",x"56",x"ED", -- 0x0650
    x"53",x"70",x"80",x"18",x"23",x"DD",x"6E",x"02", -- 0x0658
    x"DD",x"66",x"03",x"4E",x"06",x"00",x"21",x"7E", -- 0x0660
    x"0F",x"09",x"7E",x"32",x"72",x"80",x"DD",x"77", -- 0x0668
    x"01",x"18",x"0D",x"DD",x"6E",x"02",x"DD",x"66", -- 0x0670
    x"03",x"7E",x"DD",x"77",x"06",x"DD",x"77",x"07", -- 0x0678
    x"DD",x"6E",x"02",x"DD",x"66",x"03",x"23",x"DD", -- 0x0680
    x"75",x"02",x"DD",x"74",x"03",x"C3",x"09",x"0E", -- 0x0688
    x"06",x"00",x"CD",x"FE",x"05",x"DD",x"36",x"00", -- 0x0690
    x"FF",x"C9",x"CD",x"A4",x"0E",x"06",x"00",x"CD", -- 0x0698
    x"FE",x"05",x"18",x"34",x"78",x"E6",x"E0",x"07", -- 0x06A0
    x"07",x"07",x"47",x"3E",x"01",x"10",x"04",x"DD", -- 0x06A8
    x"77",x"00",x"C9",x"07",x"18",x"F7",x"C5",x"CD", -- 0x06B0
    x"A4",x"0E",x"C1",x"78",x"E6",x"1F",x"3D",x"07", -- 0x06B8
    x"4F",x"06",x"00",x"2A",x"70",x"80",x"09",x"5E", -- 0x06C0
    x"23",x"56",x"EB",x"CD",x"C6",x"04",x"DD",x"46", -- 0x06C8
    x"06",x"78",x"DD",x"77",x"07",x"CD",x"FE",x"05", -- 0x06D0
    x"DD",x"6E",x"02",x"DD",x"66",x"03",x"23",x"DD", -- 0x06D8
    x"75",x"02",x"DD",x"74",x"03",x"C9",x"06",x"0F", -- 0x06E0
    x"0A",x"0F",x"0E",x"0F",x"12",x"0F",x"16",x"0F", -- 0x06E8
    x"1A",x"0F",x"1E",x"0F",x"22",x"0F",x"26",x"0F", -- 0x06F0
    x"2A",x"0F",x"2E",x"0F",x"32",x"0F",x"36",x"0F", -- 0x06F8
    x"3A",x"0F",x"3E",x"0F",x"42",x"0F",x"6B",x"08", -- 0x0700
    x"F2",x"07",x"80",x"07",x"14",x"07",x"AE",x"06", -- 0x0708
    x"4E",x"06",x"F3",x"05",x"9E",x"05",x"4E",x"05", -- 0x0710
    x"01",x"05",x"B9",x"04",x"76",x"04",x"36",x"04", -- 0x0718
    x"F9",x"03",x"C0",x"03",x"8A",x"03",x"57",x"03", -- 0x0720
    x"27",x"03",x"FA",x"02",x"CF",x"02",x"A7",x"02", -- 0x0728
    x"81",x"02",x"5D",x"02",x"3B",x"02",x"1B",x"02", -- 0x0730
    x"FD",x"01",x"E0",x"01",x"C5",x"01",x"AC",x"01", -- 0x0738
    x"94",x"01",x"7D",x"01",x"68",x"01",x"53",x"01", -- 0x0740
    x"40",x"01",x"2E",x"01",x"1D",x"01",x"0D",x"01", -- 0x0748
    x"FE",x"00",x"F0",x"00",x"E3",x"00",x"D6",x"00", -- 0x0750
    x"CA",x"00",x"BE",x"00",x"B4",x"00",x"AA",x"00", -- 0x0758
    x"A0",x"00",x"97",x"00",x"8F",x"00",x"87",x"00", -- 0x0760
    x"7F",x"00",x"78",x"00",x"71",x"00",x"6B",x"00", -- 0x0768
    x"65",x"00",x"5F",x"00",x"5A",x"00",x"55",x"00", -- 0x0770
    x"50",x"00",x"4C",x"00",x"47",x"00",x"57",x"42", -- 0x0778
    x"34",x"2C",x"25",x"21",x"1D",x"1A",x"0C",x"0B", -- 0x0780
    x"0A",x"09",x"08",x"07",x"06",x"05",x"21",x"C1", -- 0x0788
    x"0F",x"11",x"50",x"80",x"01",x"18",x"00",x"ED", -- 0x0790
    x"B0",x"3A",x"73",x"80",x"07",x"4F",x"07",x"07", -- 0x0798
    x"91",x"4F",x"06",x"00",x"21",x"D9",x"0F",x"09", -- 0x07A0
    x"11",x"52",x"80",x"CD",x"B7",x"0F",x"11",x"5A", -- 0x07A8
    x"80",x"CD",x"B7",x"0F",x"11",x"62",x"80",x"7E", -- 0x07B0
    x"12",x"CD",x"BE",x"0F",x"7E",x"12",x"23",x"13", -- 0x07B8
    x"C9",x"01",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x07C0
    x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
    x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x07D0
    x"00",x"EB",x"0F",x"0D",x"10",x"2D",x"10",x"5F", -- 0x07D8
    x"10",x"7C",x"10",x"97",x"10",x"D5",x"10",x"EB", -- 0x07E0
    x"10",x"FF",x"10",x"1F",x"0A",x"3F",x"0D",x"5F", -- 0x07E8
    x"09",x"AC",x"80",x"6C",x"6C",x"AC",x"80",x"6C", -- 0x07F0
    x"6C",x"8C",x"88",x"8C",x"8F",x"8C",x"88",x"8C"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
