-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_PGM_45 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_PGM_45 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"00",x"2D",x"05",x"FF",x"F7",x"1F",x"04",x"3C", -- 0x0000
    x"10",x"04",x"3D",x"10",x"04",x"3C",x"10",x"04", -- 0x0008
    x"3D",x"10",x"04",x"3C",x"10",x"04",x"3D",x"10", -- 0x0010
    x"04",x"3E",x"10",x"FF",x"06",x"20",x"04",x"BC", -- 0x0018
    x"10",x"04",x"BD",x"10",x"04",x"BC",x"10",x"04", -- 0x0020
    x"BD",x"10",x"04",x"BC",x"10",x"04",x"BD",x"10", -- 0x0028
    x"04",x"BE",x"10",x"FF",x"1E",x"20",x"DD",x"21", -- 0x0030
    x"80",x"42",x"11",x"20",x"00",x"06",x"08",x"D9", -- 0x0038
    x"CD",x"49",x"20",x"D9",x"DD",x"19",x"10",x"F7", -- 0x0040
    x"C9",x"DD",x"7E",x"00",x"DD",x"B6",x"01",x"0F", -- 0x0048
    x"D0",x"DD",x"7E",x"02",x"EF",x"69",x"20",x"B2", -- 0x0050
    x"20",x"CA",x"20",x"CB",x"20",x"E5",x"20",x"E6", -- 0x0058
    x"20",x"E7",x"20",x"2A",x"21",x"47",x"21",x"48", -- 0x0060
    x"21",x"2A",x"1B",x"41",x"DD",x"75",x"18",x"DD", -- 0x0068
    x"74",x"19",x"3A",x"16",x"41",x"E6",x"0F",x"C6", -- 0x0070
    x"F8",x"DD",x"77",x"04",x"7D",x"E6",x"1F",x"07", -- 0x0078
    x"07",x"07",x"C6",x"08",x"DD",x"77",x"03",x"DD", -- 0x0080
    x"7E",x"17",x"A7",x"28",x"15",x"3D",x"28",x"08", -- 0x0088
    x"3D",x"28",x"0A",x"21",x"5B",x"21",x"18",x"0D", -- 0x0090
    x"21",x"4F",x"21",x"18",x"08",x"21",x"55",x"21", -- 0x0098
    x"18",x"03",x"21",x"49",x"21",x"DD",x"75",x"0C", -- 0x00A0
    x"DD",x"74",x"0D",x"DD",x"36",x"0E",x"00",x"DD", -- 0x00A8
    x"34",x"02",x"CD",x"63",x"1B",x"3A",x"15",x"41", -- 0x00B0
    x"A7",x"C0",x"DD",x"34",x"04",x"DD",x"7E",x"04", -- 0x00B8
    x"C6",x"14",x"FE",x"08",x"D0",x"DD",x"36",x"02", -- 0x00C0
    x"03",x"C9",x"C9",x"DD",x"6E",x"18",x"DD",x"66", -- 0x00C8
    x"19",x"3E",x"10",x"77",x"23",x"77",x"11",x"1F", -- 0x00D0
    x"00",x"19",x"77",x"23",x"77",x"AF",x"DD",x"77", -- 0x00D8
    x"00",x"DD",x"77",x"01",x"C9",x"C9",x"C9",x"DD", -- 0x00E0
    x"7E",x"17",x"3D",x"28",x"05",x"3D",x"28",x"09", -- 0x00E8
    x"18",x"23",x"21",x"76",x"21",x"3E",x"3F",x"18", -- 0x00F0
    x"21",x"DD",x"46",x"1A",x"3E",x"4F",x"05",x"28", -- 0x00F8
    x"05",x"05",x"28",x"07",x"18",x"0A",x"21",x"8B", -- 0x0100
    x"21",x"18",x"0F",x"21",x"91",x"21",x"18",x"0A", -- 0x0108
    x"21",x"85",x"21",x"18",x"05",x"21",x"67",x"21", -- 0x0110
    x"3E",x"3F",x"DD",x"75",x"0C",x"DD",x"74",x"0D", -- 0x0118
    x"DD",x"36",x"0E",x"00",x"DD",x"77",x"0F",x"DD", -- 0x0120
    x"34",x"02",x"CD",x"63",x"1B",x"DD",x"35",x"0F", -- 0x0128
    x"28",x"10",x"3A",x"15",x"41",x"A7",x"C0",x"DD", -- 0x0130
    x"34",x"04",x"DD",x"7E",x"04",x"C6",x"14",x"FE", -- 0x0138
    x"08",x"D0",x"DD",x"36",x"02",x"03",x"C9",x"C9", -- 0x0140
    x"C9",x"02",x"1C",x"10",x"FF",x"49",x"21",x"02", -- 0x0148
    x"10",x"10",x"FF",x"4F",x"21",x"02",x"33",x"10", -- 0x0150
    x"FF",x"55",x"21",x"00",x"2F",x"06",x"00",x"26", -- 0x0158
    x"06",x"00",x"1F",x"06",x"FF",x"5B",x"21",x"02", -- 0x0160
    x"38",x"10",x"02",x"39",x"10",x"02",x"3A",x"10", -- 0x0168
    x"02",x"3B",x"10",x"FF",x"67",x"21",x"02",x"38", -- 0x0170
    x"10",x"02",x"39",x"10",x"02",x"3A",x"10",x"02", -- 0x0178
    x"3B",x"10",x"FF",x"76",x"21",x"02",x"11",x"50", -- 0x0180
    x"FF",x"85",x"21",x"02",x"12",x"50",x"FF",x"8B", -- 0x0188
    x"21",x"02",x"13",x"50",x"FF",x"91",x"21",x"DD", -- 0x0190
    x"21",x"C0",x"43",x"11",x"20",x"00",x"06",x"02", -- 0x0198
    x"D9",x"CD",x"AA",x"21",x"D9",x"DD",x"19",x"10", -- 0x01A0
    x"F7",x"C9",x"DD",x"7E",x"00",x"DD",x"B6",x"01", -- 0x01A8
    x"0F",x"D0",x"DD",x"7E",x"02",x"EF",x"CA",x"21", -- 0x01B0
    x"F3",x"21",x"07",x"22",x"08",x"22",x"09",x"22", -- 0x01B8
    x"0A",x"22",x"0B",x"22",x"1F",x"22",x"35",x"22", -- 0x01C0
    x"36",x"22",x"3A",x"83",x"43",x"C6",x"04",x"DD", -- 0x01C8
    x"77",x"03",x"3A",x"84",x"43",x"C6",x"08",x"DD", -- 0x01D0
    x"77",x"04",x"21",x"37",x"22",x"DD",x"75",x"0C", -- 0x01D8
    x"DD",x"74",x"0D",x"DD",x"36",x"0E",x"00",x"21", -- 0x01E0
    x"5E",x"22",x"DD",x"75",x"13",x"DD",x"74",x"14", -- 0x01E8
    x"DD",x"34",x"02",x"CD",x"63",x"1B",x"CD",x"F7", -- 0x01F0
    x"1C",x"DD",x"7E",x"03",x"FE",x"F0",x"D8",x"AF", -- 0x01F8
    x"DD",x"77",x"00",x"DD",x"77",x"01",x"C9",x"C9", -- 0x0200
    x"C9",x"C9",x"C9",x"21",x"4F",x"22",x"DD",x"75", -- 0x0208
    x"0C",x"DD",x"74",x"0D",x"DD",x"36",x"0E",x"00", -- 0x0210
    x"DD",x"36",x"0F",x"23",x"DD",x"34",x"02",x"CD", -- 0x0218
    x"63",x"1B",x"DD",x"35",x"0F",x"20",x"05",x"AF", -- 0x0220
    x"DD",x"77",x"01",x"C9",x"3A",x"15",x"41",x"A7", -- 0x0228
    x"C0",x"DD",x"34",x"04",x"C9",x"C9",x"C9",x"06", -- 0x0230
    x"21",x"04",x"06",x"22",x"04",x"06",x"21",x"04", -- 0x0238
    x"06",x"22",x"04",x"06",x"23",x"08",x"06",x"24", -- 0x0240
    x"08",x"06",x"25",x"FE",x"FF",x"37",x"22",x"06", -- 0x0248
    x"38",x"09",x"06",x"39",x"09",x"06",x"3A",x"09", -- 0x0250
    x"06",x"3B",x"09",x"FF",x"4F",x"22",x"00",x"00", -- 0x0258
    x"01",x"00",x"00",x"FF",x"00",x"FF",x"00",x"FF", -- 0x0260
    x"00",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"FF", -- 0x0268
    x"00",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"FF", -- 0x0270
    x"00",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"FF", -- 0x0278
    x"01",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"FF", -- 0x0280
    x"01",x"FF",x"00",x"FF",x"00",x"FF",x"01",x"FF", -- 0x0288
    x"00",x"FF",x"01",x"FF",x"01",x"FF",x"00",x"FF", -- 0x0290
    x"01",x"FF",x"01",x"FF",x"01",x"FF",x"01",x"00", -- 0x0298
    x"01",x"00",x"01",x"FF",x"01",x"FF",x"01",x"00", -- 0x02A0
    x"01",x"FF",x"01",x"00",x"01",x"FF",x"01",x"00", -- 0x02A8
    x"01",x"00",x"01",x"FF",x"01",x"00",x"01",x"00", -- 0x02B0
    x"01",x"00",x"01",x"00",x"80",x"B4",x"22",x"3A", -- 0x02B8
    x"1D",x"41",x"A7",x"28",x"03",x"FE",x"08",x"C0", -- 0x02C0
    x"DD",x"21",x"00",x"44",x"11",x"20",x"00",x"06", -- 0x02C8
    x"04",x"D9",x"CD",x"DB",x"22",x"D9",x"DD",x"19", -- 0x02D0
    x"10",x"F7",x"C9",x"DD",x"7E",x"00",x"DD",x"B6", -- 0x02D8
    x"01",x"0F",x"D0",x"DD",x"7E",x"02",x"EF",x"FB", -- 0x02E0
    x"22",x"14",x"23",x"40",x"23",x"40",x"23",x"40", -- 0x02E8
    x"23",x"40",x"23",x"41",x"23",x"55",x"23",x"6B", -- 0x02F0
    x"23",x"6B",x"23",x"21",x"6C",x"23",x"DD",x"75", -- 0x02F8
    x"0C",x"DD",x"74",x"0D",x"DD",x"36",x"0E",x"00", -- 0x0300
    x"21",x"84",x"23",x"DD",x"75",x"13",x"DD",x"74", -- 0x0308
    x"14",x"DD",x"34",x"02",x"CD",x"63",x"1B",x"CD", -- 0x0310
    x"F7",x"1C",x"3A",x"17",x"41",x"DD",x"77",x"16", -- 0x0318
    x"3A",x"15",x"41",x"A7",x"20",x"03",x"DD",x"34", -- 0x0320
    x"04",x"DD",x"7E",x"04",x"FE",x"F0",x"38",x"08", -- 0x0328
    x"AF",x"DD",x"77",x"00",x"DD",x"77",x"01",x"C9", -- 0x0330
    x"DD",x"7E",x"03",x"FE",x"28",x"D0",x"18",x"F0", -- 0x0338
    x"C9",x"21",x"75",x"23",x"DD",x"75",x"0C",x"DD", -- 0x0340
    x"74",x"0D",x"DD",x"36",x"0E",x"00",x"DD",x"36", -- 0x0348
    x"0F",x"3F",x"DD",x"34",x"02",x"CD",x"63",x"1B", -- 0x0350
    x"DD",x"35",x"0F",x"20",x"05",x"AF",x"DD",x"77", -- 0x0358
    x"01",x"C9",x"3A",x"15",x"41",x"A7",x"C0",x"DD", -- 0x0360
    x"34",x"04",x"C9",x"C9",x"00",x"1D",x"10",x"00", -- 0x0368
    x"1E",x"10",x"FF",x"6C",x"23",x"06",x"38",x"05", -- 0x0370
    x"06",x"39",x"05",x"06",x"3A",x"05",x"06",x"3B", -- 0x0378
    x"05",x"FF",x"75",x"23",x"FF",x"00",x"80",x"84", -- 0x0380
    x"23",x"3A",x"1D",x"41",x"FE",x"02",x"C0",x"DD", -- 0x0388
    x"21",x"00",x"44",x"11",x"20",x"00",x"06",x"04", -- 0x0390
    x"D9",x"CD",x"A2",x"23",x"D9",x"DD",x"19",x"10", -- 0x0398
    x"F7",x"C9",x"DD",x"7E",x"00",x"DD",x"B6",x"01", -- 0x03A0
    x"0F",x"D0",x"DD",x"7E",x"02",x"EF",x"C2",x"23", -- 0x03A8
    x"DB",x"23",x"EF",x"23",x"EF",x"23",x"F0",x"23", -- 0x03B0
    x"F0",x"23",x"F1",x"23",x"05",x"24",x"1B",x"24", -- 0x03B8
    x"1B",x"24",x"21",x"1C",x"24",x"DD",x"75",x"0C", -- 0x03C0
    x"DD",x"74",x"0D",x"DD",x"36",x"0E",x"00",x"21", -- 0x03C8
    x"31",x"24",x"DD",x"75",x"13",x"DD",x"74",x"14", -- 0x03D0
    x"DD",x"34",x"02",x"CD",x"63",x"1B",x"CD",x"F7", -- 0x03D8
    x"1C",x"DD",x"7E",x"04",x"FE",x"F0",x"D8",x"AF", -- 0x03E0
    x"DD",x"77",x"00",x"DD",x"77",x"01",x"C9",x"C9", -- 0x03E8
    x"C9",x"21",x"22",x"24",x"DD",x"75",x"0C",x"DD", -- 0x03F0
    x"74",x"0D",x"DD",x"36",x"0E",x"00",x"DD",x"36", -- 0x03F8
    x"0F",x"2B",x"DD",x"34",x"02",x"CD",x"63",x"1B", -- 0x0400
    x"DD",x"35",x"0F",x"20",x"05",x"AF",x"DD",x"77", -- 0x0408
    x"01",x"C9",x"3A",x"15",x"41",x"A7",x"C0",x"DD", -- 0x0410
    x"34",x"04",x"C9",x"C9",x"05",x"1A",x"10",x"FF", -- 0x0418
    x"1C",x"24",x"04",x"38",x"0B",x"04",x"39",x"0B", -- 0x0420
    x"04",x"3A",x"0B",x"04",x"3B",x"0B",x"FF",x"22", -- 0x0428
    x"24",x"FF",x"00",x"FE",x"00",x"FE",x"00",x"FE", -- 0x0430
    x"00",x"FE",x"00",x"FE",x"00",x"FE",x"00",x"FE", -- 0x0438
    x"00",x"FE",x"00",x"FE",x"02",x"FE",x"00",x"FE", -- 0x0440
    x"02",x"FE",x"00",x"FE",x"02",x"FE",x"02",x"FE", -- 0x0448
    x"02",x"FE",x"02",x"00",x"02",x"00",x"02",x"02", -- 0x0450
    x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x0458
    x"02",x"02",x"02",x"02",x"00",x"02",x"02",x"02", -- 0x0460
    x"00",x"02",x"02",x"02",x"00",x"02",x"02",x"02", -- 0x0468
    x"00",x"02",x"00",x"02",x"00",x"02",x"00",x"02", -- 0x0470
    x"00",x"02",x"02",x"02",x"00",x"02",x"00",x"02", -- 0x0478
    x"00",x"02",x"02",x"02",x"00",x"02",x"00",x"02", -- 0x0480
    x"00",x"02",x"00",x"02",x"02",x"02",x"00",x"02", -- 0x0488
    x"02",x"02",x"00",x"02",x"00",x"02",x"02",x"02", -- 0x0490
    x"02",x"02",x"02",x"00",x"02",x"00",x"02",x"00", -- 0x0498
    x"02",x"FE",x"02",x"FE",x"02",x"FE",x"02",x"FE", -- 0x04A0
    x"02",x"FE",x"00",x"FE",x"02",x"FE",x"00",x"FE", -- 0x04A8
    x"02",x"FE",x"00",x"FE",x"02",x"FE",x"00",x"FE", -- 0x04B0
    x"02",x"FE",x"00",x"FE",x"00",x"FE",x"00",x"FE", -- 0x04B8
    x"00",x"FE",x"00",x"FE",x"00",x"80",x"31",x"24", -- 0x04C0
    x"3A",x"1D",x"41",x"FE",x"01",x"C0",x"DD",x"21", -- 0x04C8
    x"00",x"44",x"11",x"20",x"00",x"06",x"04",x"D9", -- 0x04D0
    x"CD",x"E1",x"24",x"D9",x"DD",x"19",x"10",x"F7", -- 0x04D8
    x"C9",x"DD",x"7E",x"00",x"DD",x"B6",x"01",x"0F", -- 0x04E0
    x"D0",x"DD",x"7E",x"02",x"EF",x"01",x"25",x"DB", -- 0x04E8
    x"23",x"EF",x"23",x"EF",x"23",x"F0",x"23",x"F0", -- 0x04F0
    x"23",x"F1",x"23",x"05",x"24",x"1B",x"24",x"1B", -- 0x04F8
    x"24",x"21",x"1D",x"25",x"DD",x"75",x"0C",x"DD", -- 0x0500
    x"74",x"0D",x"DD",x"36",x"0E",x"00",x"21",x"32", -- 0x0508
    x"25",x"DD",x"75",x"13",x"DD",x"74",x"14",x"DD", -- 0x0510
    x"34",x"02",x"C3",x"DB",x"23",x"00",x"35",x"05", -- 0x0518
    x"00",x"36",x"05",x"00",x"37",x"05",x"00",x"30", -- 0x0520
    x"05",x"00",x"37",x"05",x"00",x"36",x"05",x"FF", -- 0x0528
    x"1D",x"25",x"00",x"04",x"80",x"32",x"25",x"CD", -- 0x0530
    x"46",x"25",x"CD",x"5B",x"25",x"CD",x"8C",x"25", -- 0x0538
    x"CD",x"96",x"25",x"C3",x"E5",x"25",x"21",x"2A", -- 0x0540
    x"40",x"06",x"19",x"3A",x"16",x"41",x"ED",x"44", -- 0x0548
    x"4F",x"3A",x"17",x"41",x"71",x"2C",x"77",x"2C", -- 0x0550
    x"10",x"FA",x"C9",x"21",x"60",x"42",x"DD",x"21", -- 0x0558
    x"80",x"42",x"11",x"20",x"00",x"06",x"08",x"CD", -- 0x0560
    x"6F",x"25",x"DD",x"19",x"10",x"F9",x"C9",x"DD", -- 0x0568
    x"7E",x"00",x"DD",x"B6",x"01",x"0F",x"36",x"00", -- 0x0570
    x"D0",x"36",x"01",x"2C",x"DD",x"7E",x"12",x"77", -- 0x0578
    x"2C",x"DD",x"7E",x"18",x"77",x"2C",x"DD",x"7E", -- 0x0580
    x"19",x"77",x"2C",x"C9",x"DD",x"21",x"80",x"43", -- 0x0588
    x"FD",x"21",x"60",x"40",x"18",x"12",x"DD",x"21", -- 0x0590
    x"00",x"44",x"FD",x"21",x"70",x"40",x"18",x"08", -- 0x0598
    x"DD",x"21",x"80",x"44",x"FD",x"21",x"70",x"40", -- 0x05A0
    x"01",x"08",x"04",x"DD",x"7E",x"00",x"DD",x"B6", -- 0x05A8
    x"01",x"0F",x"30",x"27",x"DD",x"7E",x"16",x"FD", -- 0x05B0
    x"77",x"02",x"DD",x"7E",x"03",x"91",x"FD",x"77", -- 0x05B8
    x"03",x"DD",x"7E",x"04",x"2F",x"91",x"FD",x"77", -- 0x05C0
    x"00",x"DD",x"7E",x"12",x"FD",x"77",x"01",x"11", -- 0x05C8
    x"20",x"00",x"DD",x"19",x"1E",x"04",x"FD",x"19", -- 0x05D0
    x"10",x"D1",x"C9",x"FD",x"36",x"00",x"F8",x"FD", -- 0x05D8
    x"36",x"03",x"F8",x"18",x"EA",x"DD",x"21",x"80", -- 0x05E0
    x"40",x"FD",x"21",x"00",x"45",x"06",x"07",x"CD", -- 0x05E8
    x"FD",x"25",x"11",x"04",x"00",x"DD",x"19",x"1D", -- 0x05F0
    x"FD",x"19",x"10",x"F3",x"C9",x"FD",x"CB",x"00", -- 0x05F8
    x"46",x"28",x"23",x"FD",x"7E",x"02",x"2F",x"DD", -- 0x0600
    x"77",x"01",x"FD",x"7E",x"01",x"C6",x"05",x"DD", -- 0x0608
    x"77",x"03",x"3A",x"0F",x"40",x"0F",x"30",x"06", -- 0x0610
    x"3A",x"0D",x"40",x"0F",x"38",x"11",x"DD",x"7E", -- 0x0618
    x"03",x"2F",x"DD",x"77",x"03",x"C9",x"DD",x"36", -- 0x0620
    x"01",x"00",x"DD",x"36",x"03",x"00",x"C9",x"DD", -- 0x0628
    x"7E",x"03",x"D6",x"0D",x"DD",x"77",x"03",x"C9", -- 0x0630
    x"CD",x"60",x"26",x"CD",x"C4",x"26",x"CD",x"E0", -- 0x0638
    x"26",x"CD",x"F6",x"26",x"CD",x"15",x"27",x"CD", -- 0x0640
    x"97",x"29",x"CD",x"65",x"2A",x"CD",x"F7",x"29", -- 0x0648
    x"CD",x"8B",x"28",x"CD",x"F2",x"28",x"CD",x"2C", -- 0x0650
    x"29",x"CD",x"68",x"27",x"CD",x"CC",x"27",x"C9", -- 0x0658
    x"3A",x"80",x"43",x"0F",x"D0",x"3A",x"1D",x"41", -- 0x0660
    x"FE",x"02",x"C0",x"DD",x"21",x"00",x"44",x"11", -- 0x0668
    x"20",x"00",x"06",x"04",x"CD",x"7C",x"26",x"DD", -- 0x0670
    x"19",x"10",x"F9",x"C9",x"DD",x"CB",x"00",x"46", -- 0x0678
    x"C8",x"21",x"83",x"43",x"7E",x"DD",x"96",x"03", -- 0x0680
    x"C6",x"06",x"FE",x"0D",x"D0",x"2C",x"7E",x"C6", -- 0x0688
    x"04",x"DD",x"96",x"04",x"C6",x"0D",x"FE",x"19", -- 0x0690
    x"D0",x"DD",x"CB",x"00",x"86",x"DD",x"CB",x"01", -- 0x0698
    x"C6",x"DD",x"36",x"02",x"06",x"2D",x"2D",x"36", -- 0x06A0
    x"06",x"2D",x"36",x"01",x"2D",x"36",x"00",x"21", -- 0x06A8
    x"A0",x"43",x"36",x"00",x"2C",x"36",x"01",x"DD", -- 0x06B0
    x"36",x"17",x"00",x"3E",x"FF",x"32",x"15",x"41", -- 0x06B8
    x"CD",x"EE",x"30",x"C9",x"3A",x"80",x"43",x"0F", -- 0x06C0
    x"D0",x"3A",x"1D",x"41",x"FE",x"01",x"C0",x"DD", -- 0x06C8
    x"21",x"00",x"44",x"11",x"20",x"00",x"06",x"04", -- 0x06D0
    x"CD",x"7C",x"26",x"DD",x"19",x"10",x"F9",x"C9", -- 0x06D8
    x"3A",x"80",x"43",x"0F",x"D0",x"DD",x"21",x"80", -- 0x06E0
    x"42",x"11",x"20",x"00",x"06",x"08",x"CD",x"7C", -- 0x06E8
    x"26",x"DD",x"19",x"10",x"F9",x"C9",x"3A",x"80", -- 0x06F0
    x"43",x"0F",x"D0",x"3A",x"1D",x"41",x"A7",x"28", -- 0x06F8
    x"03",x"FE",x"08",x"C0",x"DD",x"21",x"00",x"44", -- 0x0700
    x"11",x"20",x"00",x"06",x"04",x"CD",x"7C",x"26", -- 0x0708
    x"DD",x"19",x"10",x"F9",x"C9",x"3A",x"80",x"43", -- 0x0710
    x"0F",x"D0",x"3A",x"16",x"41",x"47",x"3A",x"84", -- 0x0718
    x"43",x"D6",x"04",x"90",x"E6",x"F8",x"0F",x"0F", -- 0x0720
    x"C6",x"C0",x"6F",x"26",x"41",x"06",x"03",x"3A", -- 0x0728
    x"83",x"43",x"C6",x"03",x"5F",x"D6",x"06",x"57", -- 0x0730
    x"7E",x"BB",x"38",x"10",x"2C",x"7E",x"BA",x"30", -- 0x0738
    x"0B",x"2C",x"28",x"03",x"10",x"F2",x"C9",x"2E", -- 0x0740
    x"C0",x"10",x"ED",x"C9",x"21",x"80",x"43",x"36", -- 0x0748
    x"00",x"2C",x"36",x"01",x"2C",x"36",x"06",x"21", -- 0x0750
    x"A0",x"43",x"36",x"00",x"2C",x"36",x"01",x"3E", -- 0x0758
    x"FF",x"32",x"15",x"41",x"CD",x"EE",x"30",x"C9", -- 0x0760
    x"3A",x"1D",x"41",x"FE",x"02",x"C0",x"FD",x"21", -- 0x0768
    x"00",x"45",x"06",x"04",x"11",x"20",x"00",x"CD", -- 0x0770
    x"83",x"27",x"FD",x"23",x"FD",x"23",x"FD",x"23", -- 0x0778
    x"10",x"F5",x"C9",x"FD",x"CB",x"00",x"46",x"C8", -- 0x0780
    x"DD",x"21",x"00",x"44",x"0E",x"04",x"D9",x"CD", -- 0x0788
    x"99",x"27",x"D9",x"DD",x"19",x"0D",x"20",x"F6", -- 0x0790
    x"C9",x"DD",x"CB",x"00",x"46",x"C8",x"FD",x"7E", -- 0x0798
    x"01",x"DD",x"96",x"03",x"C6",x"03",x"FE",x"07", -- 0x07A0
    x"D0",x"FD",x"7E",x"02",x"DD",x"96",x"04",x"C6", -- 0x07A8
    x"04",x"FE",x"09",x"D0",x"DD",x"36",x"00",x"00", -- 0x07B0
    x"DD",x"36",x"01",x"01",x"DD",x"36",x"02",x"06", -- 0x07B8
    x"FD",x"36",x"00",x"00",x"11",x"08",x"03",x"FF", -- 0x07C0
    x"CD",x"E6",x"30",x"C9",x"FD",x"21",x"00",x"45", -- 0x07C8
    x"06",x"04",x"11",x"20",x"00",x"CD",x"E1",x"27", -- 0x07D0
    x"FD",x"23",x"FD",x"23",x"FD",x"23",x"10",x"F5", -- 0x07D8
    x"C9",x"FD",x"CB",x"00",x"46",x"C8",x"DD",x"21", -- 0x07E0
    x"80",x"42",x"0E",x"08",x"D9",x"CD",x"F7",x"27", -- 0x07E8
    x"D9",x"DD",x"19",x"0D",x"20",x"F6",x"C9",x"DD", -- 0x07F0
    x"CB",x"00",x"46",x"C8",x"FD",x"7E",x"01",x"DD", -- 0x07F8
    x"96",x"03",x"C6",x"07",x"FE",x"0F",x"D0",x"FD", -- 0x0800
    x"7E",x"02",x"DD",x"96",x"04",x"C6",x"04",x"FE", -- 0x0808
    x"09",x"D0",x"DD",x"36",x"00",x"00",x"DD",x"36", -- 0x0810
    x"01",x"01",x"DD",x"36",x"02",x"06",x"FD",x"36", -- 0x0818
    x"00",x"00",x"DD",x"7E",x"17",x"A7",x"28",x"08", -- 0x0820
    x"3D",x"28",x"0D",x"3D",x"28",x"1D",x"18",x"4E", -- 0x0828
    x"11",x"01",x"03",x"FF",x"CD",x"F6",x"30",x"C9", -- 0x0830
    x"21",x"05",x"41",x"7E",x"C6",x"30",x"30",x"02", -- 0x0838
    x"3E",x"FF",x"77",x"11",x"03",x"03",x"FF",x"CD", -- 0x0840
    x"C9",x"30",x"C9",x"ED",x"5F",x"E6",x"03",x"A7", -- 0x0848
    x"28",x"08",x"3D",x"28",x"05",x"3D",x"28",x"0E", -- 0x0850
    x"18",x"18",x"DD",x"36",x"1A",x"00",x"11",x"05", -- 0x0858
    x"03",x"FF",x"CD",x"D1",x"30",x"C9",x"DD",x"36", -- 0x0860
    x"1A",x"01",x"11",x"06",x"03",x"FF",x"CD",x"D1", -- 0x0868
    x"30",x"C9",x"DD",x"36",x"1A",x"02",x"11",x"07", -- 0x0870
    x"03",x"FF",x"CD",x"D1",x"30",x"C9",x"11",x"0D", -- 0x0878
    x"03",x"FF",x"CD",x"D1",x"30",x"3E",x"FF",x"32", -- 0x0880
    x"12",x"41",x"C9",x"3A",x"1D",x"41",x"A7",x"28", -- 0x0888
    x"03",x"FE",x"08",x"C0",x"FD",x"21",x"00",x"45", -- 0x0890
    x"06",x"04",x"11",x"20",x"00",x"CD",x"A9",x"28", -- 0x0898
    x"FD",x"23",x"FD",x"23",x"FD",x"23",x"10",x"F5", -- 0x08A0
    x"C9",x"FD",x"CB",x"00",x"46",x"C8",x"DD",x"21", -- 0x08A8
    x"00",x"44",x"0E",x"04",x"D9",x"CD",x"BF",x"28", -- 0x08B0
    x"D9",x"DD",x"19",x"0D",x"20",x"F6",x"C9",x"DD", -- 0x08B8
    x"CB",x"00",x"46",x"C8",x"FD",x"7E",x"01",x"DD", -- 0x08C0
    x"96",x"03",x"C6",x"05",x"FE",x"0B",x"D0",x"FD", -- 0x08C8
    x"7E",x"02",x"DD",x"96",x"04",x"C6",x"03",x"FE", -- 0x08D0
    x"07",x"D0",x"DD",x"36",x"00",x"00",x"DD",x"36", -- 0x08D8
    x"01",x"01",x"DD",x"36",x"02",x"06",x"FD",x"36", -- 0x08E0
    x"00",x"00",x"11",x"0A",x"03",x"FF",x"CD",x"F6", -- 0x08E8
    x"30",x"C9",x"DD",x"21",x"00",x"45",x"11",x"03", -- 0x08F0
    x"00",x"06",x"04",x"D9",x"CD",x"05",x"29",x"D9", -- 0x08F8
    x"DD",x"19",x"10",x"F7",x"C9",x"DD",x"CB",x"00", -- 0x0900
    x"46",x"C8",x"3A",x"16",x"41",x"47",x"DD",x"7E", -- 0x0908
    x"02",x"90",x"E6",x"F8",x"0F",x"0F",x"C6",x"C0", -- 0x0910
    x"6F",x"26",x"41",x"7E",x"DD",x"BE",x"01",x"38", -- 0x0918
    x"06",x"2C",x"7E",x"DD",x"BE",x"01",x"D8",x"DD", -- 0x0920
    x"36",x"00",x"00",x"C9",x"3A",x"1D",x"41",x"FE", -- 0x0928
    x"02",x"C0",x"FD",x"21",x"C0",x"43",x"06",x"02", -- 0x0930
    x"11",x"20",x"00",x"CD",x"43",x"29",x"FD",x"19", -- 0x0938
    x"10",x"F9",x"C9",x"FD",x"CB",x"00",x"46",x"C8", -- 0x0940
    x"DD",x"21",x"00",x"44",x"0E",x"04",x"D9",x"CD", -- 0x0948
    x"59",x"29",x"D9",x"DD",x"19",x"0D",x"20",x"F6", -- 0x0950
    x"C9",x"DD",x"CB",x"00",x"46",x"C8",x"FD",x"7E", -- 0x0958
    x"03",x"DD",x"96",x"03",x"C6",x"05",x"FE",x"0B", -- 0x0960
    x"D0",x"FD",x"7E",x"04",x"DD",x"96",x"04",x"C6", -- 0x0968
    x"06",x"FE",x"0D",x"D0",x"DD",x"36",x"00",x"00", -- 0x0970
    x"DD",x"36",x"01",x"01",x"DD",x"36",x"02",x"06", -- 0x0978
    x"FD",x"36",x"00",x"00",x"FD",x"36",x"01",x"01", -- 0x0980
    x"FD",x"36",x"02",x"06",x"11",x"08",x"03",x"FF", -- 0x0988
    x"CD",x"D9",x"30",x"CD",x"E6",x"30",x"C9",x"FD", -- 0x0990
    x"21",x"C0",x"43",x"06",x"02",x"11",x"20",x"00", -- 0x0998
    x"CD",x"A8",x"29",x"FD",x"19",x"10",x"F9",x"C9", -- 0x09A0
    x"FD",x"CB",x"00",x"46",x"C8",x"DD",x"21",x"80", -- 0x09A8
    x"42",x"0E",x"08",x"D9",x"CD",x"BE",x"29",x"D9", -- 0x09B0
    x"DD",x"19",x"0D",x"20",x"F6",x"C9",x"DD",x"CB", -- 0x09B8
    x"00",x"46",x"C8",x"FD",x"7E",x"03",x"DD",x"96", -- 0x09C0
    x"03",x"C6",x"07",x"FE",x"0E",x"D0",x"FD",x"7E", -- 0x09C8
    x"04",x"DD",x"96",x"04",x"C6",x"07",x"FE",x"0E", -- 0x09D0
    x"D0",x"DD",x"36",x"00",x"00",x"DD",x"36",x"01", -- 0x09D8
    x"01",x"DD",x"36",x"02",x"06",x"FD",x"36",x"00", -- 0x09E0
    x"00",x"FD",x"36",x"01",x"01",x"FD",x"36",x"02", -- 0x09E8
    x"06",x"CD",x"D9",x"30",x"C3",x"22",x"28",x"3A", -- 0x09F0
    x"1D",x"41",x"A7",x"28",x"03",x"FE",x"08",x"C0", -- 0x09F8
    x"FD",x"21",x"C0",x"43",x"06",x"02",x"11",x"20", -- 0x0A00
    x"00",x"CD",x"11",x"2A",x"FD",x"19",x"10",x"F9", -- 0x0A08
    x"C9",x"FD",x"CB",x"00",x"46",x"C8",x"DD",x"21", -- 0x0A10
    x"00",x"44",x"0E",x"04",x"D9",x"CD",x"27",x"2A", -- 0x0A18
    x"D9",x"DD",x"19",x"0D",x"20",x"F6",x"C9",x"DD", -- 0x0A20
    x"CB",x"00",x"46",x"C8",x"FD",x"7E",x"03",x"DD", -- 0x0A28
    x"96",x"03",x"C6",x"06",x"FE",x"0D",x"D0",x"FD", -- 0x0A30
    x"7E",x"04",x"DD",x"96",x"04",x"C6",x"04",x"FE", -- 0x0A38
    x"09",x"D0",x"DD",x"36",x"00",x"00",x"DD",x"36", -- 0x0A40
    x"01",x"01",x"DD",x"36",x"02",x"06",x"FD",x"36", -- 0x0A48
    x"00",x"00",x"FD",x"36",x"01",x"01",x"FD",x"36", -- 0x0A50
    x"02",x"06",x"11",x"0A",x"03",x"FF",x"CD",x"D9", -- 0x0A58
    x"30",x"CD",x"F6",x"30",x"C9",x"DD",x"21",x"C0", -- 0x0A60
    x"43",x"06",x"02",x"11",x"20",x"00",x"D9",x"CD", -- 0x0A68
    x"78",x"2A",x"D9",x"DD",x"19",x"10",x"F7",x"C9", -- 0x0A70
    x"DD",x"CB",x"00",x"46",x"C8",x"3A",x"16",x"41", -- 0x0A78
    x"47",x"DD",x"7E",x"04",x"90",x"E6",x"F8",x"0F", -- 0x0A80
    x"0F",x"C6",x"C0",x"6F",x"26",x"41",x"7E",x"DD", -- 0x0A88
    x"BE",x"03",x"38",x"06",x"2C",x"7E",x"DD",x"BE", -- 0x0A90
    x"03",x"D8",x"DD",x"36",x"00",x"00",x"DD",x"36", -- 0x0A98
    x"01",x"01",x"DD",x"36",x"02",x"06",x"CD",x"D9", -- 0x0AA0
    x"30",x"C9",x"3A",x"06",x"40",x"0F",x"38",x"19", -- 0x0AA8
    x"3A",x"80",x"43",x"0F",x"30",x"19",x"3A",x"5F", -- 0x0AB0
    x"42",x"E6",x"67",x"CC",x"0A",x"2B",x"3A",x"5F", -- 0x0AB8
    x"42",x"E6",x"3F",x"CC",x"38",x"2C",x"C3",x"CF", -- 0x0AC0
    x"2A",x"CD",x"13",x"2C",x"CD",x"E5",x"2A",x"CD", -- 0x0AC8
    x"2D",x"2B",x"CD",x"6A",x"2B",x"CD",x"D6",x"2B", -- 0x0AD0
    x"CD",x"57",x"2C",x"CD",x"5C",x"2F",x"CD",x"2A", -- 0x0AD8
    x"2F",x"CD",x"8E",x"2F",x"C9",x"3A",x"80",x"43", -- 0x0AE0
    x"0F",x"D0",x"3A",x"0D",x"40",x"0F",x"38",x"0E", -- 0x0AE8
    x"3A",x"10",x"40",x"CB",x"5F",x"C8",x"3A",x"13", -- 0x0AF0
    x"40",x"CB",x"5F",x"C0",x"18",x"0C",x"3A",x"11", -- 0x0AF8
    x"40",x"CB",x"5F",x"C8",x"3A",x"14",x"40",x"CB", -- 0x0B00
    x"5F",x"C0",x"21",x"00",x"45",x"06",x"04",x"CB", -- 0x0B08
    x"46",x"20",x"14",x"CB",x"C6",x"2C",x"3A",x"83", -- 0x0B10
    x"43",x"C6",x"02",x"77",x"2C",x"3A",x"84",x"43", -- 0x0B18
    x"D6",x"07",x"77",x"CD",x"FE",x"30",x"C9",x"2C", -- 0x0B20
    x"2C",x"2C",x"10",x"E3",x"C9",x"3A",x"1D",x"41", -- 0x0B28
    x"FE",x"02",x"C0",x"3A",x"5F",x"42",x"E6",x"3F", -- 0x0B30
    x"C0",x"DD",x"21",x"00",x"44",x"11",x"20",x"00", -- 0x0B38
    x"06",x"04",x"DD",x"7E",x"00",x"DD",x"B6",x"01", -- 0x0B40
    x"0F",x"30",x"05",x"DD",x"19",x"10",x"F3",x"C9", -- 0x0B48
    x"DD",x"36",x"00",x"01",x"DD",x"36",x"01",x"00", -- 0x0B50
    x"DD",x"36",x"02",x"00",x"DD",x"36",x"03",x"88", -- 0x0B58
    x"ED",x"5F",x"E6",x"0F",x"C6",x"09",x"DD",x"77", -- 0x0B60
    x"04",x"C9",x"3A",x"1D",x"41",x"A7",x"28",x"03", -- 0x0B68
    x"FE",x"08",x"C0",x"3A",x"5F",x"42",x"E6",x"1F", -- 0x0B70
    x"C0",x"ED",x"5F",x"E6",x"01",x"C8",x"DD",x"21", -- 0x0B78
    x"80",x"42",x"11",x"20",x"00",x"06",x"08",x"DD", -- 0x0B80
    x"CB",x"00",x"46",x"20",x"05",x"DD",x"19",x"10", -- 0x0B88
    x"F6",x"C9",x"DD",x"7E",x"17",x"A7",x"20",x"F5", -- 0x0B90
    x"3A",x"A4",x"43",x"DD",x"96",x"04",x"FE",x"70", -- 0x0B98
    x"30",x"EB",x"FD",x"21",x"00",x"44",x"06",x"04", -- 0x0BA0
    x"FD",x"7E",x"00",x"FD",x"B6",x"01",x"0F",x"30", -- 0x0BA8
    x"05",x"FD",x"19",x"10",x"F3",x"C9",x"DD",x"36", -- 0x0BB0
    x"02",x"03",x"DD",x"7E",x"03",x"FD",x"77",x"03", -- 0x0BB8
    x"DD",x"7E",x"04",x"FD",x"77",x"04",x"FD",x"36", -- 0x0BC0
    x"00",x"01",x"FD",x"36",x"01",x"00",x"FD",x"36", -- 0x0BC8
    x"02",x"00",x"CD",x"08",x"31",x"C9",x"3A",x"1D", -- 0x0BD0
    x"41",x"FE",x"01",x"C0",x"3A",x"5F",x"42",x"E6", -- 0x0BD8
    x"0F",x"C0",x"DD",x"21",x"00",x"44",x"11",x"20", -- 0x0BE0
    x"00",x"06",x"04",x"DD",x"7E",x"00",x"DD",x"B6", -- 0x0BE8
    x"01",x"0F",x"30",x"05",x"DD",x"19",x"10",x"F3", -- 0x0BF0
    x"C9",x"DD",x"36",x"00",x"01",x"DD",x"36",x"01", -- 0x0BF8
    x"00",x"DD",x"36",x"02",x"00",x"ED",x"5F",x"E6", -- 0x0C00
    x"7F",x"C6",x"30",x"DD",x"77",x"03",x"DD",x"36", -- 0x0C08
    x"04",x"08",x"C9",x"3A",x"80",x"43",x"0F",x"D0", -- 0x0C10
    x"3A",x"0D",x"40",x"0F",x"38",x"0E",x"3A",x"10", -- 0x0C18
    x"40",x"CB",x"4F",x"C8",x"3A",x"13",x"40",x"CB", -- 0x0C20
    x"4F",x"C0",x"18",x"0C",x"3A",x"11",x"40",x"CB", -- 0x0C28
    x"57",x"C8",x"3A",x"14",x"40",x"CB",x"57",x"C0", -- 0x0C30
    x"21",x"C0",x"43",x"11",x"1F",x"00",x"06",x"02", -- 0x0C38
    x"7E",x"2C",x"B6",x"0F",x"30",x"04",x"19",x"10", -- 0x0C40
    x"F7",x"C9",x"2D",x"36",x"01",x"2C",x"36",x"00", -- 0x0C48
    x"2C",x"36",x"00",x"CD",x"03",x"31",x"C9",x"3A", -- 0x0C50
    x"1A",x"41",x"E6",x"02",x"C8",x"DD",x"21",x"80", -- 0x0C58
    x"42",x"11",x"20",x"00",x"06",x"08",x"DD",x"7E", -- 0x0C60
    x"00",x"DD",x"B6",x"01",x"0F",x"30",x"05",x"DD", -- 0x0C68
    x"19",x"10",x"F3",x"C9",x"DD",x"36",x"00",x"01", -- 0x0C70
    x"DD",x"36",x"01",x"00",x"DD",x"36",x"02",x"00", -- 0x0C78
    x"DD",x"36",x"17",x"01",x"AF",x"32",x"1A",x"41", -- 0x0C80
    x"C9",x"C8",x"36",x"CB",x"2E",x"00",x"00",x"D3", -- 0x0C88
    x"2C",x"DB",x"2E",x"00",x"00",x"E0",x"36",x"E0", -- 0x0C90
    x"36",x"00",x"01",x"DB",x"30",x"D3",x"33",x"00", -- 0x0C98
    x"00",x"D0",x"35",x"CB",x"32",x"00",x"00",x"C3", -- 0x0CA0
    x"33",x"B8",x"30",x"00",x"00",x"BB",x"2F",x"C3", -- 0x0CA8
    x"2D",x"00",x"00",x"CB",x"2E",x"D3",x"2C",x"00", -- 0x0CB0
    x"00",x"DB",x"2E",x"E0",x"36",x"00",x"00",x"E0", -- 0x0CB8
    x"36",x"E0",x"36",x"00",x"01",x"E0",x"36",x"E0", -- 0x0CC0
    x"36",x"00",x"02",x"E0",x"36",x"E0",x"36",x"00", -- 0x0CC8
    x"01",x"DB",x"30",x"D0",x"32",x"00",x"00",x"D3", -- 0x0CD0
    x"2E",x"DB",x"2C",x"00",x"00",x"DB",x"30",x"D3", -- 0x0CD8
    x"32",x"00",x"00",x"C8",x"34",x"D3",x"2F",x"00", -- 0x0CE0
    x"00",x"D8",x"36",x"D8",x"36",x"00",x"02",x"D3", -- 0x0CE8
    x"30",x"CB",x"33",x"00",x"00",x"C3",x"30",x"BB", -- 0x0CF0
    x"33",x"00",x"00",x"B8",x"2F",x"B8",x"30",x"00", -- 0x0CF8
    x"00",x"B8",x"2E",x"C3",x"2D",x"00",x"00",x"CB", -- 0x0D00
    x"2C",x"D3",x"2F",x"00",x"00",x"D8",x"36",x"D8", -- 0x0D08
    x"36",x"00",x"01",x"D8",x"36",x"DB",x"2E",x"00", -- 0x0D10
    x"00",x"E0",x"36",x"E0",x"36",x"00",x"04",x"E0", -- 0x0D18
    x"36",x"E0",x"36",x"00",x"02",x"E0",x"36",x"DB", -- 0x0D20
    x"33",x"00",x"00",x"D3",x"30",x"C8",x"30",x"00", -- 0x0D28
    x"00",x"C0",x"33",x"B8",x"34",x"00",x"00",x"C3", -- 0x0D30
    x"2F",x"CB",x"2D",x"00",x"00",x"D3",x"2C",x"DB", -- 0x0D38
    x"2F",x"00",x"00",x"E0",x"36",x"E0",x"36",x"00", -- 0x0D40
    x"02",x"D8",x"32",x"D8",x"35",x"00",x"00",x"DB", -- 0x0D48
    x"2C",x"E0",x"36",x"00",x"00",x"E0",x"36",x"E0", -- 0x0D50
    x"36",x"00",x"04",x"E0",x"36",x"E0",x"36",x"00", -- 0x0D58
    x"04",x"E0",x"36",x"D8",x"34",x"00",x"00",x"E0", -- 0x0D60
    x"36",x"E0",x"36",x"00",x"02",x"E0",x"36",x"E0", -- 0x0D68
    x"36",x"00",x"01",x"E0",x"36",x"E0",x"36",x"00", -- 0x0D70
    x"01",x"D8",x"32",x"D8",x"35",x"00",x"00",x"D0", -- 0x0D78
    x"30",x"D0",x"2D",x"00",x"00",x"DB",x"2F",x"E0", -- 0x0D80
    x"36",x"00",x"00",x"E0",x"36",x"E0",x"36",x"00", -- 0x0D88
    x"04",x"E0",x"36",x"E0",x"36",x"00",x"04",x"E0", -- 0x0D90
    x"36",x"E0",x"36",x"00",x"01",x"E0",x"36",x"E0", -- 0x0D98
    x"36",x"00",x"02",x"E0",x"36",x"E0",x"36",x"00", -- 0x0DA0
    x"01",x"DB",x"30",x"D3",x"31",x"00",x"00",x"CB", -- 0x0DA8
    x"32",x"C3",x"33",x"00",x"00",x"BB",x"31",x"BB", -- 0x0DB0
    x"2C",x"00",x"00",x"C3",x"2D",x"CB",x"2E",x"00", -- 0x0DB8
    x"00",x"D0",x"2C",x"D8",x"2E",x"00",x"00",x"E0", -- 0x0DC0
    x"36",x"E0",x"36",x"00",x"02",x"E0",x"36",x"DB", -- 0x0DC8
    x"33",x"00",x"00",x"D0",x"33",x"CB",x"33",x"00", -- 0x0DD0
    x"00",x"C8",x"36",x"CB",x"2E",x"00",x"00",x"D3", -- 0x0DD8
    x"2C",x"DB",x"2E",x"00",x"00",x"E0",x"36",x"E0", -- 0x0DE0
    x"36",x"00",x"04",x"DB",x"30",x"D3",x"33",x"00", -- 0x0DE8
    x"00",x"D0",x"35",x"CB",x"32",x"00",x"00",x"C3", -- 0x0DF0
    x"33",x"B8",x"30",x"00",x"00",x"BB",x"2F",x"C3", -- 0x0DF8
    x"2D",x"00",x"00",x"CB",x"2E",x"D3",x"2C",x"00", -- 0x0E00
    x"00",x"DB",x"2E",x"E0",x"36",x"00",x"00",x"E0", -- 0x0E08
    x"36",x"E0",x"36",x"00",x"02",x"E0",x"36",x"E0", -- 0x0E10
    x"36",x"00",x"01",x"E0",x"36",x"E0",x"36",x"00", -- 0x0E18
    x"01",x"DB",x"30",x"D0",x"32",x"00",x"00",x"D3", -- 0x0E20
    x"2E",x"DB",x"2C",x"00",x"00",x"DB",x"30",x"D3", -- 0x0E28
    x"32",x"00",x"00",x"C8",x"34",x"D3",x"2F",x"00", -- 0x0E30
    x"00",x"D8",x"36",x"D8",x"36",x"00",x"02",x"D3", -- 0x0E38
    x"30",x"CB",x"33",x"00",x"00",x"C3",x"30",x"BB", -- 0x0E40
    x"33",x"00",x"00",x"B8",x"2F",x"B8",x"30",x"00", -- 0x0E48
    x"00",x"B8",x"2E",x"C3",x"2D",x"00",x"00",x"CB", -- 0x0E50
    x"2C",x"D3",x"2F",x"00",x"00",x"D8",x"36",x"D8", -- 0x0E58
    x"36",x"00",x"00",x"D8",x"36",x"DB",x"2E",x"00", -- 0x0E60
    x"00",x"E0",x"36",x"E0",x"36",x"00",x"04",x"E0", -- 0x0E68
    x"36",x"E0",x"36",x"00",x"02",x"E0",x"36",x"DB", -- 0x0E70
    x"33",x"00",x"00",x"D3",x"30",x"C8",x"30",x"00", -- 0x0E78
    x"00",x"C8",x"36",x"CB",x"2E",x"00",x"00",x"D3", -- 0x0E80
    x"2C",x"DB",x"2E",x"00",x"00",x"E0",x"36",x"E0", -- 0x0E88
    x"36",x"00",x"01",x"DB",x"30",x"D3",x"33",x"00", -- 0x0E90
    x"00",x"D0",x"35",x"CB",x"32",x"00",x"00",x"C3", -- 0x0E98
    x"33",x"B8",x"30",x"00",x"00",x"BB",x"2F",x"C3", -- 0x0EA0
    x"2D",x"00",x"00",x"CB",x"2E",x"D3",x"2C",x"00", -- 0x0EA8
    x"00",x"DB",x"2E",x"E0",x"36",x"00",x"00",x"E0", -- 0x0EB0
    x"36",x"E0",x"36",x"00",x"01",x"E0",x"36",x"E0", -- 0x0EB8
    x"36",x"00",x"01",x"E0",x"36",x"E0",x"36",x"00", -- 0x0EC0
    x"02",x"DB",x"30",x"D0",x"32",x"00",x"00",x"D3", -- 0x0EC8
    x"2E",x"DB",x"2C",x"00",x"00",x"DB",x"30",x"D3", -- 0x0ED0
    x"32",x"00",x"00",x"C8",x"34",x"D3",x"2F",x"00", -- 0x0ED8
    x"00",x"D8",x"36",x"D8",x"36",x"00",x"02",x"D3", -- 0x0EE0
    x"30",x"CB",x"33",x"00",x"00",x"C3",x"30",x"BB", -- 0x0EE8
    x"33",x"00",x"00",x"B8",x"2F",x"B8",x"30",x"00", -- 0x0EF0
    x"00",x"B8",x"2E",x"C3",x"2D",x"00",x"00",x"CB", -- 0x0EF8
    x"2C",x"D3",x"2F",x"00",x"00",x"D8",x"36",x"D8", -- 0x0F00
    x"36",x"00",x"00",x"D8",x"36",x"DB",x"2E",x"00", -- 0x0F08
    x"00",x"E0",x"36",x"E0",x"36",x"00",x"02",x"E0", -- 0x0F10
    x"36",x"E0",x"36",x"00",x"04",x"E0",x"36",x"DB", -- 0x0F18
    x"33",x"00",x"00",x"D3",x"30",x"C8",x"30",x"00", -- 0x0F20
    x"00",x"FF",x"3A",x"1A",x"41",x"E6",x"01",x"C8", -- 0x0F28
    x"DD",x"21",x"80",x"42",x"11",x"20",x"00",x"06", -- 0x0F30
    x"08",x"DD",x"7E",x"00",x"DD",x"B6",x"01",x"0F", -- 0x0F38
    x"30",x"05",x"DD",x"19",x"10",x"F3",x"C9",x"DD", -- 0x0F40
    x"36",x"00",x"01",x"DD",x"36",x"01",x"00",x"DD", -- 0x0F48
    x"36",x"02",x"00",x"DD",x"36",x"17",x"00",x"AF", -- 0x0F50
    x"32",x"1A",x"41",x"C9",x"3A",x"1A",x"41",x"E6", -- 0x0F58
    x"04",x"C8",x"DD",x"21",x"80",x"42",x"11",x"20", -- 0x0F60
    x"00",x"06",x"08",x"DD",x"7E",x"00",x"DD",x"B6", -- 0x0F68
    x"01",x"0F",x"30",x"05",x"DD",x"19",x"10",x"F3", -- 0x0F70
    x"C9",x"DD",x"36",x"00",x"01",x"DD",x"36",x"01", -- 0x0F78
    x"00",x"DD",x"36",x"02",x"00",x"DD",x"36",x"17", -- 0x0F80
    x"02",x"AF",x"32",x"1A",x"41",x"C9",x"3A",x"1A", -- 0x0F88
    x"41",x"E6",x"08",x"C8",x"DD",x"21",x"80",x"42", -- 0x0F90
    x"11",x"20",x"00",x"06",x"08",x"DD",x"7E",x"00", -- 0x0F98
    x"DD",x"B6",x"01",x"0F",x"30",x"05",x"DD",x"19", -- 0x0FA0
    x"10",x"F3",x"C9",x"DD",x"36",x"00",x"01",x"DD", -- 0x0FA8
    x"36",x"01",x"00",x"DD",x"36",x"02",x"00",x"DD", -- 0x0FB0
    x"36",x"17",x"03",x"AF",x"32",x"1A",x"41",x"C9", -- 0x0FB8
    x"CD",x"C7",x"2F",x"CD",x"02",x"30",x"C9",x"2A", -- 0x0FC0
    x"18",x"41",x"7E",x"FE",x"FF",x"C0",x"21",x"00", -- 0x0FC8
    x"44",x"11",x"01",x"44",x"01",x"80",x"00",x"36", -- 0x0FD0
    x"00",x"ED",x"B0",x"21",x"1E",x"41",x"7E",x"FE", -- 0x0FD8
    x"05",x"28",x"01",x"34",x"7E",x"47",x"87",x"80", -- 0x0FE0
    x"5F",x"16",x"00",x"21",x"B5",x"31",x"19",x"7E", -- 0x0FE8
    x"32",x"18",x"41",x"23",x"7E",x"32",x"19",x"41", -- 0x0FF0
    x"23",x"7E",x"32",x"1D",x"41",x"11",x"02",x"07"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
