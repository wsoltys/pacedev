-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_PGM_67 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_PGM_67 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"FF",x"C9",x"3A",x"5F",x"42",x"A7",x"C0",x"21", -- 0x0000
    x"1B",x"40",x"34",x"7E",x"0F",x"D8",x"21",x"17", -- 0x0008
    x"41",x"7E",x"3C",x"E6",x"07",x"FE",x"01",x"28", -- 0x0010
    x"03",x"77",x"18",x"02",x"3C",x"77",x"47",x"3A", -- 0x0018
    x"11",x"41",x"0F",x"38",x"13",x"78",x"21",x"40", -- 0x0020
    x"30",x"16",x"00",x"87",x"5F",x"19",x"7E",x"32", -- 0x0028
    x"04",x"68",x"23",x"7E",x"32",x"03",x"68",x"C9", -- 0x0030
    x"AF",x"32",x"04",x"68",x"32",x"03",x"68",x"C9", -- 0x0038
    x"01",x"00",x"01",x"00",x"01",x"00",x"01",x"00", -- 0x0040
    x"01",x"01",x"01",x"01",x"01",x"00",x"01",x"00", -- 0x0048
    x"11",x"41",x"42",x"1A",x"6F",x"26",x"42",x"7E", -- 0x0050
    x"FE",x"FF",x"C8",x"47",x"3A",x"06",x"40",x"A7", -- 0x0058
    x"78",x"C4",x"AD",x"30",x"36",x"FF",x"7D",x"FE", -- 0x0060
    x"5E",x"28",x"03",x"3C",x"12",x"C9",x"3E",x"43", -- 0x0068
    x"12",x"C9",x"C5",x"D5",x"E5",x"47",x"11",x"40", -- 0x0070
    x"42",x"1A",x"6F",x"26",x"42",x"70",x"7D",x"FE", -- 0x0078
    x"5E",x"28",x"04",x"3C",x"12",x"18",x"03",x"3E", -- 0x0080
    x"43",x"12",x"E1",x"D1",x"C1",x"C9",x"3A",x"42", -- 0x0088
    x"42",x"F6",x"10",x"32",x"42",x"42",x"32",x"01", -- 0x0090
    x"82",x"AF",x"C3",x"AD",x"30",x"AF",x"CD",x"AD", -- 0x0098
    x"30",x"3A",x"42",x"42",x"E6",x"EF",x"32",x"42", -- 0x00A0
    x"42",x"32",x"01",x"82",x"C9",x"32",x"00",x"82", -- 0x00A8
    x"3A",x"42",x"42",x"E6",x"F7",x"32",x"01",x"82", -- 0x00B0
    x"00",x"00",x"00",x"00",x"3A",x"42",x"42",x"F6", -- 0x00B8
    x"08",x"32",x"01",x"82",x"C9",x"3E",x"08",x"18", -- 0x00C0
    x"E4",x"3E",x"01",x"CD",x"72",x"30",x"C3",x"31", -- 0x00C8
    x"31",x"3E",x"01",x"CD",x"72",x"30",x"C3",x"31", -- 0x00D0
    x"31",x"3E",x"30",x"CD",x"72",x"30",x"3E",x"02", -- 0x00D8
    x"CD",x"72",x"30",x"C3",x"31",x"31",x"3E",x"04", -- 0x00E0
    x"CD",x"72",x"30",x"C3",x"31",x"31",x"3E",x"05", -- 0x00E8
    x"CD",x"72",x"30",x"C3",x"31",x"31",x"3E",x"03", -- 0x00F0
    x"CD",x"72",x"30",x"C3",x"31",x"31",x"3E",x"06", -- 0x00F8
    x"C3",x"72",x"30",x"3E",x"20",x"C3",x"72",x"30", -- 0x0100
    x"C9",x"3E",x"0A",x"C3",x"72",x"30",x"3E",x"09", -- 0x0108
    x"CD",x"72",x"30",x"3E",x"0A",x"C3",x"72",x"30", -- 0x0110
    x"3E",x"0B",x"CD",x"72",x"30",x"3E",x"0C",x"CD", -- 0x0118
    x"72",x"30",x"3E",x"0D",x"C3",x"72",x"30",x"3E", -- 0x0120
    x"0E",x"CD",x"72",x"30",x"3E",x"0F",x"C3",x"72", -- 0x0128
    x"30",x"3E",x"13",x"CD",x"72",x"30",x"3E",x"14", -- 0x0130
    x"CD",x"72",x"30",x"3E",x"15",x"C3",x"72",x"30", -- 0x0138
    x"3A",x"42",x"42",x"F6",x"40",x"B0",x"32",x"42", -- 0x0140
    x"42",x"32",x"01",x"82",x"C9",x"3A",x"42",x"42", -- 0x0148
    x"E6",x"BF",x"32",x"42",x"42",x"32",x"01",x"82", -- 0x0150
    x"AF",x"32",x"1C",x"40",x"C9",x"3E",x"12",x"C3", -- 0x0158
    x"72",x"30",x"3E",x"21",x"C3",x"72",x"30",x"3E", -- 0x0160
    x"07",x"C3",x"72",x"30",x"3E",x"22",x"CD",x"72", -- 0x0168
    x"30",x"3E",x"23",x"C3",x"72",x"30",x"3E",x"24", -- 0x0170
    x"C3",x"72",x"30",x"3A",x"5F",x"42",x"E6",x"3F", -- 0x0178
    x"C0",x"3A",x"05",x"41",x"FE",x"50",x"DC",x"67", -- 0x0180
    x"31",x"3A",x"1D",x"41",x"FE",x"00",x"CC",x"5D", -- 0x0188
    x"31",x"FE",x"01",x"CC",x"6C",x"31",x"FE",x"02", -- 0x0190
    x"28",x"0D",x"FE",x"04",x"CC",x"76",x"31",x"FE", -- 0x0198
    x"08",x"CC",x"5D",x"31",x"C3",x"5D",x"31",x"3A", -- 0x01A0
    x"5F",x"42",x"E6",x"7F",x"CA",x"62",x"31",x"C9", -- 0x01A8
    x"3E",x"08",x"C3",x"72",x"30",x"C7",x"31",x"00", -- 0x01B0
    x"0E",x"14",x"02",x"89",x"2C",x"01",x"ED",x"06", -- 0x01B8
    x"08",x"B8",x"35",x"04",x"A9",x"39",x"10",x"C0", -- 0x01C0
    x"33",x"BC",x"31",x"00",x"00",x"B0",x"32",x"AB", -- 0x01C8
    x"31",x"00",x"00",x"A0",x"33",x"9B",x"30",x"00", -- 0x01D0
    x"00",x"93",x"30",x"8B",x"33",x"00",x"00",x"83", -- 0x01D8
    x"30",x"7B",x"31",x"00",x"00",x"70",x"32",x"68", -- 0x01E0
    x"32",x"00",x"00",x"60",x"34",x"6B",x"2D",x"00", -- 0x01E8
    x"00",x"73",x"2D",x"7B",x"2E",x"00",x"00",x"80", -- 0x01F0
    x"36",x"80",x"36",x"00",x"01",x"83",x"2C",x"83", -- 0x01F8
    x"30",x"00",x"00",x"80",x"36",x"80",x"36",x"00", -- 0x0200
    x"01",x"80",x"36",x"80",x"36",x"00",x"00",x"80", -- 0x0208
    x"36",x"80",x"36",x"00",x"01",x"80",x"36",x"80", -- 0x0210
    x"36",x"00",x"00",x"80",x"36",x"80",x"36",x"00", -- 0x0218
    x"01",x"80",x"36",x"80",x"36",x"00",x"01",x"80", -- 0x0220
    x"36",x"80",x"36",x"00",x"01",x"80",x"35",x"80", -- 0x0228
    x"35",x"00",x"00",x"80",x"36",x"80",x"36",x"00", -- 0x0230
    x"02",x"83",x"35",x"7B",x"30",x"00",x"00",x"73", -- 0x0238
    x"30",x"6B",x"31",x"00",x"00",x"60",x"32",x"60", -- 0x0240
    x"2C",x"00",x"00",x"6B",x"2C",x"73",x"2C",x"00", -- 0x0248
    x"00",x"7B",x"2F",x"83",x"2F",x"00",x"00",x"8B", -- 0x0250
    x"2E",x"93",x"2D",x"00",x"00",x"98",x"2E",x"A0", -- 0x0258
    x"2E",x"00",x"00",x"AB",x"2D",x"B0",x"2F",x"00", -- 0x0260
    x"00",x"BB",x"2C",x"C3",x"2C",x"00",x"00",x"C8", -- 0x0268
    x"36",x"C8",x"2E",x"00",x"00",x"D3",x"2D",x"DB", -- 0x0270
    x"2E",x"00",x"00",x"E0",x"36",x"E0",x"36",x"00", -- 0x0278
    x"01",x"E0",x"36",x"E0",x"36",x"00",x"01",x"D8", -- 0x0280
    x"32",x"D8",x"35",x"00",x"00",x"DB",x"2C",x"E0", -- 0x0288
    x"36",x"00",x"00",x"E0",x"36",x"E0",x"36",x"00", -- 0x0290
    x"02",x"E0",x"36",x"E0",x"36",x"00",x"02",x"E0", -- 0x0298
    x"36",x"D8",x"34",x"00",x"00",x"E0",x"36",x"E0", -- 0x02A0
    x"36",x"00",x"01",x"E0",x"36",x"E0",x"36",x"00", -- 0x02A8
    x"01",x"E0",x"36",x"E0",x"36",x"00",x"04",x"D8", -- 0x02B0
    x"32",x"D8",x"35",x"00",x"00",x"D0",x"30",x"D0", -- 0x02B8
    x"2D",x"00",x"00",x"DB",x"2F",x"E0",x"36",x"00", -- 0x02C0
    x"00",x"E0",x"36",x"E0",x"36",x"00",x"00",x"E0", -- 0x02C8
    x"36",x"E0",x"36",x"00",x"01",x"E0",x"36",x"E0", -- 0x02D0
    x"36",x"00",x"00",x"E0",x"36",x"E0",x"36",x"00", -- 0x02D8
    x"01",x"E0",x"36",x"E0",x"36",x"00",x"00",x"E0", -- 0x02E0
    x"36",x"E0",x"36",x"00",x"01",x"E0",x"36",x"E0", -- 0x02E8
    x"36",x"00",x"04",x"E0",x"36",x"E0",x"36",x"00", -- 0x02F0
    x"02",x"D8",x"30",x"D3",x"30",x"00",x"00",x"D0", -- 0x02F8
    x"2C",x"D8",x"2E",x"00",x"00",x"E0",x"36",x"E0", -- 0x0300
    x"36",x"00",x"01",x"E0",x"36",x"DB",x"33",x"00", -- 0x0308
    x"00",x"D0",x"33",x"CB",x"33",x"00",x"00",x"C8", -- 0x0310
    x"36",x"C8",x"36",x"00",x"01",x"C0",x"31",x"C0", -- 0x0318
    x"36",x"00",x"00",x"C0",x"36",x"C0",x"36",x"00", -- 0x0320
    x"01",x"B9",x"34",x"C0",x"35",x"00",x"00",x"C0", -- 0x0328
    x"36",x"C0",x"36",x"00",x"01",x"B8",x"34",x"B8", -- 0x0330
    x"33",x"00",x"00",x"B8",x"36",x"B8",x"36",x"00", -- 0x0338
    x"01",x"B8",x"36",x"B8",x"36",x"00",x"01",x"B0", -- 0x0340
    x"33",x"A8",x"34",x"00",x"00",x"B0",x"36",x"B0", -- 0x0348
    x"36",x"00",x"04",x"B0",x"36",x"B0",x"36",x"00", -- 0x0350
    x"02",x"A8",x"33",x"A0",x"32",x"00",x"00",x"A0", -- 0x0358
    x"36",x"A0",x"36",x"00",x"01",x"A0",x"36",x"A0", -- 0x0360
    x"36",x"00",x"01",x"98",x"34",x"98",x"30",x"00", -- 0x0368
    x"00",x"98",x"2C",x"98",x"33",x"00",x"00",x"98", -- 0x0370
    x"36",x"98",x"36",x"00",x"01",x"98",x"36",x"98", -- 0x0378
    x"36",x"00",x"01",x"90",x"34",x"90",x"33",x"00", -- 0x0380
    x"00",x"90",x"36",x"90",x"36",x"00",x"01",x"90", -- 0x0388
    x"36",x"90",x"36",x"00",x"01",x"8B",x"32",x"83", -- 0x0390
    x"31",x"00",x"00",x"7B",x"33",x"73",x"34",x"00", -- 0x0398
    x"00",x"7B",x"2D",x"83",x"2E",x"00",x"00",x"8B", -- 0x03A0
    x"2D",x"93",x"2F",x"00",x"00",x"9B",x"2C",x"A3", -- 0x03A8
    x"2E",x"00",x"00",x"AB",x"2C",x"B3",x"2D",x"00", -- 0x03B0
    x"00",x"B8",x"36",x"B8",x"36",x"00",x"01",x"B8", -- 0x03B8
    x"36",x"B8",x"36",x"00",x"01",x"B3",x"32",x"AB", -- 0x03C0
    x"33",x"00",x"00",x"A0",x"34",x"A0",x"34",x"00", -- 0x03C8
    x"00",x"A8",x"36",x"A8",x"36",x"00",x"01",x"A3", -- 0x03D0
    x"32",x"9B",x"32",x"00",x"00",x"90",x"34",x"98", -- 0x03D8
    x"35",x"00",x"00",x"98",x"36",x"98",x"36",x"00", -- 0x03E0
    x"01",x"93",x"30",x"8B",x"33",x"00",x"00",x"83", -- 0x03E8
    x"32",x"7B",x"30",x"00",x"00",x"73",x"33",x"6B", -- 0x03F0
    x"31",x"00",x"00",x"60",x"34",x"6B",x"2E",x"00", -- 0x03F8
    x"00",x"70",x"35",x"70",x"2E",x"00",x"00",x"78", -- 0x0400
    x"36",x"78",x"36",x"00",x"01",x"7B",x"2D",x"83", -- 0x0408
    x"2D",x"00",x"00",x"88",x"36",x"88",x"36",x"00", -- 0x0410
    x"02",x"8B",x"2F",x"93",x"2D",x"00",x"00",x"9B", -- 0x0418
    x"2E",x"A0",x"35",x"00",x"00",x"A0",x"36",x"A0", -- 0x0420
    x"36",x"00",x"01",x"A3",x"2C",x"A3",x"30",x"00", -- 0x0428
    x"00",x"9B",x"33",x"90",x"33",x"00",x"00",x"90", -- 0x0430
    x"36",x"90",x"36",x"00",x"01",x"90",x"36",x"90", -- 0x0438
    x"36",x"00",x"04",x"88",x"30",x"88",x"2C",x"00", -- 0x0440
    x"00",x"90",x"36",x"90",x"36",x"00",x"01",x"88", -- 0x0448
    x"34",x"93",x"2E",x"00",x"00",x"9B",x"2D",x"A3", -- 0x0450
    x"2F",x"00",x"00",x"AB",x"2C",x"B3",x"2E",x"00", -- 0x0458
    x"00",x"BB",x"2F",x"C3",x"2C",x"00",x"00",x"C8", -- 0x0460
    x"36",x"CB",x"2E",x"00",x"00",x"D0",x"36",x"D0", -- 0x0468
    x"36",x"00",x"01",x"D0",x"35",x"C8",x"34",x"00", -- 0x0470
    x"00",x"D0",x"36",x"D0",x"36",x"00",x"02",x"D0", -- 0x0478
    x"36",x"D0",x"36",x"00",x"02",x"CB",x"31",x"C3", -- 0x0480
    x"33",x"00",x"00",x"C0",x"36",x"C0",x"36",x"00", -- 0x0488
    x"01",x"C0",x"36",x"BB",x"32",x"00",x"00",x"B0", -- 0x0490
    x"30",x"B0",x"2E",x"00",x"00",x"B8",x"36",x"B3", -- 0x0498
    x"33",x"00",x"00",x"AB",x"32",x"AB",x"2C",x"00", -- 0x04A0
    x"00",x"B3",x"2C",x"BB",x"2C",x"00",x"00",x"C3", -- 0x04A8
    x"2C",x"C8",x"36",x"00",x"00",x"C8",x"36",x"C8", -- 0x04B0
    x"36",x"00",x"01",x"C8",x"36",x"C8",x"35",x"00", -- 0x04B8
    x"00",x"C8",x"36",x"C0",x"34",x"00",x"00",x"CB", -- 0x04C0
    x"2C",x"D3",x"2C",x"00",x"00",x"DB",x"2C",x"DB", -- 0x04C8
    x"30",x"00",x"00",x"D8",x"36",x"D8",x"36",x"00", -- 0x04D0
    x"02",x"DB",x"2D",x"E0",x"36",x"00",x"00",x"E0", -- 0x04D8
    x"36",x"E0",x"36",x"00",x"04",x"D8",x"34",x"D8", -- 0x04E0
    x"30",x"00",x"00",x"D8",x"36",x"D8",x"36",x"00", -- 0x04E8
    x"01",x"D3",x"30",x"CB",x"32",x"00",x"00",x"C8", -- 0x04F0
    x"36",x"C8",x"36",x"00",x"01",x"C8",x"36",x"C8", -- 0x04F8
    x"36",x"00",x"04",x"CB",x"2C",x"D0",x"35",x"00", -- 0x0500
    x"00",x"CB",x"30",x"C8",x"36",x"00",x"00",x"C0", -- 0x0508
    x"33",x"BB",x"33",x"00",x"00",x"B3",x"31",x"AB", -- 0x0510
    x"33",x"00",x"00",x"A0",x"34",x"A8",x"35",x"00", -- 0x0518
    x"00",x"A8",x"36",x"A8",x"36",x"00",x"01",x"A8", -- 0x0520
    x"36",x"A8",x"36",x"00",x"01",x"A8",x"36",x"A8", -- 0x0528
    x"36",x"00",x"04",x"A8",x"36",x"A8",x"36",x"00", -- 0x0530
    x"02",x"A8",x"35",x"A8",x"2C",x"00",x"00",x"B0", -- 0x0538
    x"36",x"B0",x"36",x"00",x"01",x"B0",x"36",x"B0", -- 0x0540
    x"36",x"00",x"01",x"B0",x"36",x"B0",x"36",x"00", -- 0x0548
    x"01",x"B0",x"36",x"B0",x"36",x"00",x"00",x"A8", -- 0x0550
    x"34",x"A8",x"31",x"00",x"00",x"A8",x"36",x"A8", -- 0x0558
    x"36",x"00",x"02",x"A8",x"36",x"A8",x"36",x"00", -- 0x0560
    x"01",x"A8",x"36",x"A8",x"36",x"00",x"04",x"AB", -- 0x0568
    x"2F",x"B3",x"2E",x"00",x"00",x"BB",x"2D",x"C0", -- 0x0570
    x"35",x"00",x"00",x"C0",x"36",x"C0",x"36",x"00", -- 0x0578
    x"02",x"BB",x"31",x"B3",x"32",x"00",x"00",x"AB", -- 0x0580
    x"31",x"A0",x"34",x"00",x"00",x"A3",x"31",x"9B", -- 0x0588
    x"32",x"00",x"00",x"93",x"33",x"90",x"35",x"00", -- 0x0590
    x"00",x"8B",x"32",x"80",x"34",x"00",x"00",x"8B", -- 0x0598
    x"2C",x"93",x"2E",x"00",x"00",x"9B",x"2F",x"A3", -- 0x05A0
    x"2C",x"00",x"00",x"AB",x"2D",x"B3",x"2E",x"00", -- 0x05A8
    x"00",x"BB",x"2D",x"C3",x"2F",x"00",x"00",x"FF", -- 0x05B0
    x"60",x"D1",x"60",x"D1",x"47",x"D1",x"47",x"D1", -- 0x05B8
    x"02",x"60",x"D1",x"60",x"D1",x"47",x"D1",x"47", -- 0x05C0
    x"D1",x"02",x"60",x"D1",x"60",x"D1",x"37",x"D1", -- 0x05C8
    x"37",x"D1",x"00",x"60",x"D1",x"60",x"D1",x"37", -- 0x05D0
    x"D1",x"37",x"D1",x"00",x"60",x"D1",x"60",x"D1", -- 0x05D8
    x"37",x"D1",x"37",x"D1",x"00",x"50",x"D1",x"50", -- 0x05E0
    x"D1",x"37",x"D1",x"37",x"D1",x"02",x"50",x"D1", -- 0x05E8
    x"50",x"D1",x"37",x"D1",x"37",x"D1",x"00",x"60", -- 0x05F0
    x"D1",x"60",x"D1",x"37",x"D1",x"37",x"D1",x"00", -- 0x05F8
    x"60",x"D1",x"60",x"D1",x"37",x"D1",x"37",x"D1", -- 0x0600
    x"00",x"60",x"D1",x"60",x"D1",x"37",x"D1",x"37", -- 0x0608
    x"D1",x"00",x"60",x"D1",x"60",x"D1",x"47",x"D1", -- 0x0610
    x"47",x"D1",x"00",x"60",x"D1",x"60",x"D1",x"47", -- 0x0618
    x"D1",x"47",x"D1",x"00",x"60",x"D1",x"60",x"D1", -- 0x0620
    x"47",x"D1",x"47",x"D1",x"02",x"60",x"D1",x"60", -- 0x0628
    x"D1",x"47",x"D1",x"47",x"D1",x"02",x"60",x"D1", -- 0x0630
    x"60",x"D1",x"47",x"D1",x"47",x"D1",x"02",x"60", -- 0x0638
    x"D1",x"60",x"D1",x"2F",x"D1",x"2F",x"D1",x"02", -- 0x0640
    x"60",x"D1",x"60",x"D1",x"2F",x"D1",x"2F",x"D1", -- 0x0648
    x"00",x"60",x"D1",x"60",x"D1",x"2F",x"D1",x"2F", -- 0x0650
    x"D1",x"00",x"40",x"D1",x"40",x"D1",x"2F",x"D1", -- 0x0658
    x"2F",x"D1",x"00",x"40",x"D1",x"40",x"D1",x"2F", -- 0x0660
    x"D1",x"2F",x"D1",x"00",x"40",x"D1",x"40",x"D1", -- 0x0668
    x"2F",x"D1",x"2F",x"D1",x"00",x"40",x"D1",x"40", -- 0x0670
    x"D1",x"2F",x"D1",x"2F",x"D1",x"00",x"40",x"D1", -- 0x0678
    x"40",x"D1",x"2F",x"D1",x"2F",x"D1",x"00",x"A0", -- 0x0680
    x"D1",x"A0",x"D1",x"2F",x"D1",x"2F",x"D1",x"00", -- 0x0688
    x"A0",x"D1",x"A0",x"D1",x"2F",x"D1",x"2F",x"D1", -- 0x0690
    x"00",x"A0",x"D1",x"A0",x"D1",x"2F",x"D1",x"2F", -- 0x0698
    x"D1",x"00",x"A0",x"D1",x"A0",x"D1",x"2F",x"D1", -- 0x06A0
    x"2F",x"D1",x"00",x"A0",x"D1",x"A0",x"D1",x"2F", -- 0x06A8
    x"D1",x"2F",x"D1",x"02",x"A0",x"D1",x"A0",x"D1", -- 0x06B0
    x"2F",x"D1",x"2F",x"D1",x"02",x"A0",x"D1",x"A0", -- 0x06B8
    x"D1",x"37",x"D1",x"37",x"D1",x"02",x"A0",x"D1", -- 0x06C0
    x"A0",x"D1",x"8F",x"D1",x"8F",x"D1",x"02",x"A0", -- 0x06C8
    x"D1",x"A0",x"D1",x"8F",x"D1",x"8F",x"D1",x"02", -- 0x06D0
    x"A0",x"D1",x"A0",x"D1",x"8F",x"D1",x"8F",x"D1", -- 0x06D8
    x"02",x"A0",x"D1",x"A0",x"D1",x"8F",x"D1",x"8F", -- 0x06E0
    x"D1",x"00",x"A0",x"D1",x"A0",x"D1",x"8F",x"D1", -- 0x06E8
    x"8F",x"D1",x"00",x"A0",x"D1",x"A0",x"D1",x"8F", -- 0x06F0
    x"D1",x"8F",x"D1",x"00",x"D8",x"D1",x"D8",x"D1", -- 0x06F8
    x"8F",x"D1",x"8F",x"D1",x"00",x"D8",x"D1",x"D8", -- 0x0700
    x"D1",x"8F",x"D1",x"8F",x"D1",x"00",x"D8",x"D1", -- 0x0708
    x"D8",x"D1",x"8F",x"D1",x"8F",x"D1",x"00",x"D8", -- 0x0710
    x"D1",x"D8",x"D1",x"C7",x"D1",x"C7",x"D1",x"00", -- 0x0718
    x"D8",x"D1",x"D8",x"D1",x"C7",x"D1",x"C7",x"D1", -- 0x0720
    x"02",x"D8",x"D1",x"D8",x"D1",x"C7",x"D1",x"C7", -- 0x0728
    x"D1",x"02",x"D8",x"D1",x"D8",x"D1",x"C7",x"D1", -- 0x0730
    x"C7",x"D1",x"02",x"D8",x"D1",x"D8",x"D1",x"C7", -- 0x0738
    x"D1",x"C7",x"D1",x"02",x"D8",x"D1",x"D8",x"D1", -- 0x0740
    x"C7",x"D1",x"C7",x"D1",x"00",x"D8",x"D1",x"D8", -- 0x0748
    x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"D8",x"D1", -- 0x0750
    x"D8",x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"D8", -- 0x0758
    x"D1",x"D8",x"D1",x"3F",x"D1",x"3F",x"D1",x"00", -- 0x0760
    x"D8",x"D1",x"D8",x"D1",x"3F",x"D1",x"3F",x"D1", -- 0x0768
    x"00",x"D8",x"D1",x"D8",x"D1",x"3F",x"D1",x"3F", -- 0x0770
    x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"3F",x"D1", -- 0x0778
    x"3F",x"D1",x"00",x"50",x"D1",x"50",x"D1",x"3F", -- 0x0780
    x"D1",x"3F",x"D1",x"00",x"50",x"D1",x"50",x"D1", -- 0x0788
    x"3F",x"D1",x"3F",x"D1",x"00",x"50",x"D1",x"50", -- 0x0790
    x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"50",x"D1", -- 0x0798
    x"50",x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"50", -- 0x07A0
    x"D1",x"50",x"D1",x"3F",x"D1",x"3F",x"D1",x"00", -- 0x07A8
    x"D8",x"D1",x"D8",x"D1",x"3F",x"D1",x"3F",x"D1", -- 0x07B0
    x"00",x"D8",x"D1",x"D8",x"D1",x"3F",x"D1",x"3F", -- 0x07B8
    x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"3F",x"D1", -- 0x07C0
    x"3F",x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"3F", -- 0x07C8
    x"D1",x"3F",x"D1",x"00",x"D8",x"D1",x"D8",x"D1", -- 0x07D0
    x"3F",x"D1",x"3F",x"D1",x"00",x"D8",x"D1",x"D8", -- 0x07D8
    x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"D8",x"D1", -- 0x07E0
    x"D8",x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"D8", -- 0x07E8
    x"D1",x"D8",x"D1",x"C7",x"D1",x"C7",x"D1",x"00", -- 0x07F0
    x"D8",x"D1",x"D8",x"D1",x"C7",x"D1",x"C7",x"D1", -- 0x07F8
    x"00",x"D8",x"D1",x"D8",x"D1",x"C7",x"D1",x"C7", -- 0x0800
    x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"C7",x"D1", -- 0x0808
    x"C7",x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"C7", -- 0x0810
    x"D1",x"C7",x"D1",x"00",x"D8",x"D1",x"D8",x"D1", -- 0x0818
    x"C7",x"D1",x"C7",x"D1",x"00",x"D8",x"D1",x"D8", -- 0x0820
    x"D1",x"C7",x"D1",x"C7",x"D1",x"00",x"D8",x"D1", -- 0x0828
    x"D8",x"D1",x"4F",x"D1",x"4F",x"D1",x"00",x"D8", -- 0x0830
    x"D1",x"D8",x"D1",x"4F",x"D1",x"4F",x"D1",x"00", -- 0x0838
    x"D8",x"D1",x"D8",x"D1",x"4F",x"D1",x"4F",x"D1", -- 0x0840
    x"00",x"D8",x"D1",x"D8",x"D1",x"4F",x"D1",x"4F", -- 0x0848
    x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"4F",x"D1", -- 0x0850
    x"4F",x"D1",x"00",x"60",x"D1",x"60",x"D1",x"4F", -- 0x0858
    x"D1",x"4F",x"D1",x"00",x"60",x"D1",x"60",x"D1", -- 0x0860
    x"4F",x"D1",x"4F",x"D1",x"00",x"60",x"D1",x"60", -- 0x0868
    x"D1",x"4F",x"D1",x"4F",x"D1",x"00",x"60",x"D1", -- 0x0870
    x"60",x"D1",x"37",x"D1",x"37",x"D1",x"00",x"60", -- 0x0878
    x"D1",x"60",x"D1",x"37",x"D1",x"37",x"D1",x"00", -- 0x0880
    x"48",x"D1",x"48",x"D1",x"37",x"D1",x"37",x"D1", -- 0x0888
    x"00",x"48",x"D1",x"48",x"D1",x"37",x"D1",x"37", -- 0x0890
    x"D1",x"00",x"48",x"D1",x"48",x"D1",x"37",x"D1", -- 0x0898
    x"37",x"D1",x"00",x"58",x"D1",x"58",x"D1",x"37", -- 0x08A0
    x"D1",x"37",x"D1",x"00",x"58",x"D1",x"58",x"D1", -- 0x08A8
    x"37",x"D1",x"37",x"D1",x"00",x"58",x"D1",x"58", -- 0x08B0
    x"D1",x"47",x"D1",x"47",x"D1",x"00",x"58",x"D1", -- 0x08B8
    x"58",x"D1",x"47",x"D1",x"47",x"D1",x"00",x"58", -- 0x08C0
    x"D1",x"58",x"D1",x"47",x"D1",x"47",x"D1",x"00", -- 0x08C8
    x"58",x"D1",x"58",x"D1",x"47",x"D1",x"47",x"D1", -- 0x08D0
    x"00",x"D8",x"D1",x"D8",x"D1",x"47",x"D1",x"47", -- 0x08D8
    x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"47",x"D1", -- 0x08E0
    x"47",x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"47", -- 0x08E8
    x"D1",x"47",x"D1",x"00",x"D8",x"D1",x"D8",x"D1", -- 0x08F0
    x"47",x"D1",x"47",x"D1",x"00",x"D8",x"D1",x"D8", -- 0x08F8
    x"D1",x"47",x"D1",x"47",x"D1",x"00",x"D8",x"D1", -- 0x0900
    x"D8",x"D1",x"C7",x"D1",x"C7",x"D1",x"00",x"D8", -- 0x0908
    x"D1",x"D8",x"D1",x"C7",x"D1",x"C7",x"D1",x"00", -- 0x0910
    x"D8",x"D1",x"D8",x"D1",x"C7",x"D1",x"C7",x"D1", -- 0x0918
    x"00",x"D8",x"D1",x"D8",x"D1",x"C7",x"D1",x"C7", -- 0x0920
    x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"C7",x"D1", -- 0x0928
    x"C7",x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"C7", -- 0x0930
    x"D1",x"C7",x"D1",x"02",x"D8",x"D1",x"D8",x"D1", -- 0x0938
    x"C7",x"D1",x"C7",x"D1",x"02",x"D8",x"D1",x"D8", -- 0x0940
    x"D1",x"C7",x"D1",x"C7",x"D1",x"02",x"D8",x"D1", -- 0x0948
    x"D8",x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"D8", -- 0x0950
    x"D1",x"D8",x"D1",x"3F",x"D1",x"3F",x"D1",x"00", -- 0x0958
    x"D8",x"D1",x"D8",x"D1",x"3F",x"D1",x"3F",x"D1", -- 0x0960
    x"00",x"D8",x"D1",x"D8",x"D1",x"3F",x"D1",x"3F", -- 0x0968
    x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"3F",x"D1", -- 0x0970
    x"3F",x"D1",x"00",x"D8",x"D1",x"D8",x"D1",x"3F", -- 0x0978
    x"D1",x"3F",x"D1",x"00",x"50",x"D1",x"50",x"D1", -- 0x0980
    x"3F",x"D1",x"3F",x"D1",x"00",x"60",x"D1",x"60", -- 0x0988
    x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"60",x"D1", -- 0x0990
    x"60",x"D1",x"3F",x"D1",x"3F",x"D1",x"00",x"60", -- 0x0998
    x"D1",x"60",x"D1",x"3F",x"D1",x"3F",x"D1",x"00", -- 0x09A0
    x"FF",x"C8",x"D1",x"C8",x"D1",x"00",x"00",x"C8", -- 0x09A8
    x"D1",x"C8",x"D1",x"00",x"00",x"90",x"D1",x"90", -- 0x09B0
    x"D1",x"00",x"00",x"50",x"D1",x"50",x"D1",x"00", -- 0x09B8
    x"00",x"90",x"D1",x"90",x"D1",x"00",x"00",x"C8", -- 0x09C0
    x"D1",x"C8",x"D1",x"00",x"00",x"C8",x"D1",x"C8", -- 0x09C8
    x"D1",x"00",x"00",x"98",x"D1",x"98",x"D1",x"00", -- 0x09D0
    x"00",x"98",x"D1",x"98",x"D1",x"00",x"00",x"98", -- 0x09D8
    x"D1",x"98",x"D1",x"00",x"00",x"C8",x"D1",x"C8", -- 0x09E0
    x"D1",x"00",x"00",x"48",x"D1",x"48",x"D1",x"00", -- 0x09E8
    x"00",x"48",x"D1",x"48",x"D1",x"00",x"00",x"48", -- 0x09F0
    x"D1",x"48",x"D1",x"00",x"00",x"C8",x"D1",x"C8", -- 0x09F8
    x"D1",x"00",x"00",x"98",x"D1",x"98",x"D1",x"00", -- 0x0A00
    x"00",x"98",x"D1",x"98",x"D1",x"00",x"00",x"98", -- 0x0A08
    x"D1",x"98",x"D1",x"00",x"00",x"C8",x"D1",x"C8", -- 0x0A10
    x"D1",x"00",x"00",x"C8",x"D1",x"C8",x"D1",x"00", -- 0x0A18
    x"00",x"C8",x"D1",x"C8",x"D1",x"00",x"08",x"C8", -- 0x0A20
    x"D1",x"C8",x"D1",x"00",x"00",x"C8",x"D1",x"C8", -- 0x0A28
    x"D1",x"00",x"00",x"C8",x"D1",x"C8",x"D1",x"00", -- 0x0A30
    x"00",x"70",x"D1",x"70",x"D1",x"00",x"00",x"70", -- 0x0A38
    x"D1",x"70",x"D1",x"00",x"00",x"C8",x"D1",x"C8", -- 0x0A40
    x"D1",x"00",x"00",x"C8",x"D1",x"C8",x"D1",x"00", -- 0x0A48
    x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0ED0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
