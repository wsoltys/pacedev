-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_SND_2 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_SND_2 is


  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"88",x"91",x"8D",x"92",x"8A",x"92",x"8D",x"92", -- 0x0000
    x"8A",x"92",x"8D",x"91",x"88",x"91",x"8D",x"91", -- 0x0008
    x"88",x"91",x"8F",x"94",x"FF",x"E7",x"AF",x"32", -- 0x0010
    x"C8",x"42",x"3E",x"19",x"32",x"A3",x"42",x"F7", -- 0x0018
    x"C3",x"61",x"09",x"E7",x"F7",x"C9",x"DD",x"21", -- 0x0020
    x"80",x"42",x"C3",x"A1",x"07",x"DD",x"21",x"88", -- 0x0028
    x"42",x"C3",x"A1",x"07",x"1F",x"0B",x"3F",x"0C", -- 0x0030
    x"5F",x"05",x"B4",x"91",x"8D",x"B9",x"98",x"96", -- 0x0038
    x"B4",x"99",x"91",x"8F",x"B4",x"80",x"80",x"94", -- 0x0040
    x"94",x"94",x"94",x"91",x"8F",x"8D",x"80",x"99", -- 0x0048
    x"99",x"99",x"9B",x"99",x"98",x"96",x"94",x"91", -- 0x0050
    x"80",x"91",x"B9",x"B1",x"94",x"CF",x"80",x"A0", -- 0x0058
    x"80",x"91",x"91",x"92",x"94",x"96",x"98",x"D6", -- 0x0060
    x"C0",x"80",x"92",x"92",x"94",x"B6",x"98",x"99", -- 0x0068
    x"D8",x"A0",x"B4",x"D9",x"99",x"98",x"96",x"94", -- 0x0070
    x"D8",x"B6",x"B6",x"B4",x"BB",x"B9",x"B8",x"D9", -- 0x0078
    x"C0",x"99",x"99",x"99",x"99",x"99",x"99",x"98", -- 0x0080
    x"96",x"D9",x"B4",x"91",x"91",x"AF",x"8F",x"8F", -- 0x0088
    x"99",x"99",x"98",x"96",x"D6",x"D4",x"94",x"91", -- 0x0090
    x"91",x"91",x"B1",x"8F",x"8D",x"92",x"91",x"92", -- 0x0098
    x"94",x"B6",x"A0",x"94",x"92",x"8F",x"8F",x"AF", -- 0x00A0
    x"8D",x"8C",x"8D",x"8C",x"8D",x"8F",x"D1",x"94", -- 0x00A8
    x"91",x"91",x"91",x"B1",x"8F",x"8D",x"92",x"91", -- 0x00B0
    x"92",x"94",x"B6",x"98",x"96",x"B4",x"94",x"96", -- 0x00B8
    x"94",x"92",x"91",x"8F",x"CA",x"AC",x"AF",x"CD", -- 0x00C0
    x"C0",x"FF",x"1F",x"05",x"5F",x"05",x"D9",x"D6", -- 0x00C8
    x"D9",x"D8",x"8D",x"91",x"88",x"91",x"8D",x"91", -- 0x00D0
    x"88",x"91",x"8D",x"92",x"8A",x"92",x"8D",x"92", -- 0x00D8
    x"8A",x"92",x"8D",x"91",x"88",x"91",x"8D",x"91", -- 0x00E0
    x"88",x"91",x"8F",x"94",x"88",x"94",x"8A",x"94", -- 0x00E8
    x"8C",x"94",x"8D",x"91",x"88",x"91",x"8D",x"91", -- 0x00F0
    x"88",x"91",x"8D",x"92",x"8A",x"92",x"8D",x"92", -- 0x00F8
    x"8A",x"92",x"8D",x"92",x"8A",x"92",x"8D",x"92", -- 0x0100
    x"8A",x"92",x"8F",x"94",x"88",x"94",x"8F",x"94", -- 0x0108
    x"88",x"94",x"8D",x"91",x"88",x"91",x"8D",x"91", -- 0x0110
    x"88",x"91",x"8D",x"91",x"89",x"91",x"8A",x"92", -- 0x0118
    x"8F",x"92",x"8F",x"94",x"88",x"94",x"8F",x"94", -- 0x0120
    x"88",x"94",x"8D",x"91",x"88",x"91",x"AD",x"A0", -- 0x0128
    x"D2",x"C0",x"D1",x"C0",x"DF",x"C0",x"D2",x"D2", -- 0x0130
    x"8D",x"91",x"88",x"91",x"8D",x"91",x"88",x"91", -- 0x0138
    x"8D",x"92",x"8A",x"92",x"8D",x"92",x"8A",x"92", -- 0x0140
    x"8F",x"94",x"88",x"94",x"8F",x"94",x"88",x"94", -- 0x0148
    x"8D",x"91",x"88",x"91",x"8D",x"91",x"88",x"91", -- 0x0150
    x"8D",x"91",x"88",x"91",x"8D",x"91",x"88",x"91", -- 0x0158
    x"8D",x"92",x"8A",x"92",x"8D",x"92",x"8A",x"92", -- 0x0160
    x"8F",x"94",x"88",x"94",x"8F",x"94",x"88",x"94", -- 0x0168
    x"D2",x"D4",x"8D",x"FF",x"1F",x"0B",x"3F",x"0D", -- 0x0170
    x"5F",x"06",x"8F",x"60",x"6F",x"8F",x"60",x"6F", -- 0x0178
    x"91",x"60",x"71",x"93",x"60",x"73",x"74",x"74", -- 0x0180
    x"74",x"60",x"94",x"60",x"76",x"D8",x"B9",x"B9", -- 0x0188
    x"98",x"60",x"B9",x"60",x"8F",x"60",x"6F",x"91", -- 0x0190
    x"60",x"D2",x"60",x"94",x"60",x"76",x"94",x"60", -- 0x0198
    x"72",x"91",x"60",x"71",x"92",x"60",x"D4",x"60", -- 0x01A0
    x"A0",x"74",x"76",x"78",x"60",x"B9",x"B9",x"98", -- 0x01A8
    x"60",x"B9",x"60",x"8F",x"60",x"6F",x"91",x"60", -- 0x01B0
    x"72",x"80",x"60",x"76",x"94",x"60",x"73",x"94", -- 0x01B8
    x"80",x"B2",x"B1",x"8F",x"60",x"CD",x"FF",x"1F", -- 0x01C0
    x"05",x"5F",x"06",x"B9",x"B9",x"B9",x"B9",x"B8", -- 0x01C8
    x"B2",x"B1",x"AF",x"AD",x"B4",x"B6",x"B6",x"B6", -- 0x01D0
    x"B6",x"B6",x"B6",x"B8",x"B8",x"B8",x"B8",x"B4", -- 0x01D8
    x"B1",x"BD",x"B4",x"B4",x"B4",x"B6",x"B6",x"B6", -- 0x01E0
    x"B6",x"B6",x"B6",x"98",x"80",x"A0",x"B6",x"B4", -- 0x01E8
    x"FF",x"1F",x"0B",x"3F",x"0D",x"5F",x"06",x"92", -- 0x01F0
    x"97",x"97",x"99",x"9B",x"97",x"9B",x"99",x"92", -- 0x01F8
    x"97",x"97",x"99",x"9B",x"B7",x"96",x"92",x"97", -- 0x0200
    x"97",x"99",x"9B",x"9C",x"9B",x"99",x"97",x"96", -- 0x0208
    x"92",x"94",x"96",x"B7",x"97",x"80",x"FF",x"FF", -- 0x0210
    x"1F",x"0B",x"3F",x"0D",x"5F",x"06",x"94",x"60", -- 0x0218
    x"76",x"94",x"92",x"94",x"96",x"B7",x"92",x"60", -- 0x0220
    x"74",x"92",x"90",x"8F",x"90",x"92",x"80",x"94", -- 0x0228
    x"60",x"76",x"94",x"92",x"94",x"96",x"97",x"94", -- 0x0230
    x"94",x"97",x"96",x"99",x"B7",x"97",x"80",x"FF", -- 0x0238
    x"1F",x"0B",x"5F",x"06",x"90",x"60",x"70",x"90", -- 0x0240
    x"92",x"90",x"90",x"B0",x"8F",x"60",x"70",x"8F", -- 0x0248
    x"8D",x"8B",x"8B",x"8B",x"80",x"90",x"60",x"70", -- 0x0250
    x"90",x"92",x"90",x"90",x"90",x"90",x"8F",x"92", -- 0x0258
    x"92",x"90",x"AF",x"8F",x"80",x"FF",x"1F",x"0B", -- 0x0260
    x"3F",x"0D",x"5F",x"06",x"72",x"74",x"B6",x"96", -- 0x0268
    x"B6",x"96",x"B7",x"96",x"B6",x"7B",x"7B",x"B9", -- 0x0270
    x"96",x"96",x"94",x"92",x"B4",x"94",x"B4",x"80", -- 0x0278
    x"B6",x"96",x"B6",x"96",x"B7",x"96",x"B6",x"9B", -- 0x0280
    x"B9",x"96",x"94",x"96",x"94",x"B2",x"92",x"B2", -- 0x0288
    x"80",x"FF",x"1F",x"0B",x"5F",x"06",x"72",x"74", -- 0x0290
    x"B6",x"8D",x"8D",x"8F",x"8D",x"AF",x"92",x"B2", -- 0x0298
    x"80",x"AD",x"8D",x"8F",x"91",x"92",x"B2",x"91", -- 0x02A0
    x"B1",x"72",x"74",x"B6",x"8D",x"8D",x"8F",x"8D", -- 0x02A8
    x"AF",x"92",x"B2",x"97",x"B6",x"92",x"91",x"92", -- 0x02B0
    x"9D",x"AA",x"8A",x"AA",x"80",x"FF",x"1F",x"0B", -- 0x02B8
    x"3F",x"0D",x"5F",x"06",x"8A",x"AF",x"8E",x"8C", -- 0x02C0
    x"AA",x"80",x"8A",x"AC",x"AE",x"AF",x"8A",x"8A", -- 0x02C8
    x"8C",x"8A",x"88",x"87",x"8C",x"8A",x"88",x"87", -- 0x02D0
    x"A5",x"AA",x"AA",x"80",x"FF",x"1F",x"0B",x"5F", -- 0x02D8
    x"06",x"8A",x"AF",x"8E",x"8C",x"AA",x"80",x"8A", -- 0x02E0
    x"A9",x"A8",x"A7",x"87",x"83",x"88",x"87",x"85", -- 0x02E8
    x"83",x"A3",x"A5",x"A1",x"80",x"FF",x"1F",x"0B", -- 0x02F0
    x"3F",x"0D",x"5F",x"06",x"8A",x"87",x"8A",x"8A", -- 0x02F8
    x"8A",x"8C",x"8A",x"8A",x"8A",x"87",x"8A",x"8A", -- 0x0300
    x"8A",x"8C",x"8A",x"8A",x"8A",x"AF",x"B1",x"93", -- 0x0308
    x"60",x"6F",x"8F",x"8F",x"B1",x"AE",x"AF",x"80", -- 0x0310
    x"FF",x"1F",x"0B",x"5F",x"06",x"87",x"83",x"87", -- 0x0318
    x"87",x"87",x"86",x"87",x"87",x"87",x"83",x"87", -- 0x0320
    x"87",x"87",x"87",x"85",x"87",x"88",x"AA",x"AA", -- 0x0328
    x"8A",x"60",x"67",x"87",x"8A",x"A8",x"A8",x"A7", -- 0x0330
    x"80",x"FF",x"1F",x"0B",x"3F",x"0D",x"5F",x"06", -- 0x0338
    x"8F",x"93",x"B6",x"B6",x"BB",x"9A",x"98",x"96", -- 0x0340
    x"96",x"93",x"94",x"96",x"80",x"BA",x"98",x"98", -- 0x0348
    x"94",x"98",x"96",x"96",x"9B",x"9B",x"9A",x"98", -- 0x0350
    x"96",x"9A",x"9B",x"80",x"8F",x"93",x"B6",x"B6", -- 0x0358
    x"BB",x"9A",x"98",x"96",x"96",x"93",x"94",x"96", -- 0x0360
    x"80",x"BA",x"98",x"98",x"94",x"98",x"96",x"96", -- 0x0368
    x"9B",x"9B",x"9A",x"98",x"96",x"9A",x"9B",x"80", -- 0x0370
    x"A0",x"FF",x"1F",x"0B",x"5F",x"06",x"8F",x"8F", -- 0x0378
    x"B3",x"B3",x"B8",x"96",x"94",x"93",x"93",x"8F", -- 0x0380
    x"91",x"93",x"80",x"B6",x"94",x"94",x"8F",x"94", -- 0x0388
    x"93",x"93",x"93",x"93",x"96",x"93",x"8F",x"91", -- 0x0390
    x"93",x"80",x"8F",x"8F",x"B3",x"B3",x"B8",x"96", -- 0x0398
    x"94",x"93",x"93",x"8F",x"91",x"93",x"80",x"B6", -- 0x03A0
    x"94",x"94",x"8F",x"94",x"93",x"93",x"93",x"93", -- 0x03A8
    x"96",x"93",x"8F",x"91",x"93",x"80",x"A0",x"FF", -- 0x03B0
    x"1F",x"0B",x"3F",x"0D",x"5F",x"06",x"8D",x"92", -- 0x03B8
    x"96",x"B9",x"99",x"96",x"B7",x"97",x"94",x"B6", -- 0x03C0
    x"B9",x"80",x"96",x"97",x"99",x"BB",x"9B",x"9B", -- 0x03C8
    x"9B",x"99",x"9B",x"9C",x"DD",x"A0",x"9D",x"9D", -- 0x03D0
    x"BD",x"9B",x"99",x"BB",x"99",x"97",x"9B",x"80", -- 0x03D8
    x"B9",x"A0",x"96",x"97",x"B9",x"98",x"99",x"BB", -- 0x03E0
    x"99",x"97",x"D6",x"FF",x"1F",x"0B",x"5F",x"06", -- 0x03E8
    x"8D",x"92",x"96",x"B6",x"96",x"92",x"B4",x"94", -- 0x03F0
    x"91",x"B2",x"B6",x"80",x"92",x"94",x"96",x"B7", -- 0x03F8
    x"97",x"97",x"97",x"96",x"97",x"98",x"D9",x"A0", -- 0x0400
    x"99",x"99",x"B9",x"97",x"96",x"B7",x"96",x"94", -- 0x0408
    x"97",x"80",x"B6",x"A0",x"92",x"94",x"B6",x"95", -- 0x0410
    x"96",x"B7",x"96",x"94",x"D2",x"FF",x"1F",x"0B", -- 0x0418
    x"3F",x"0D",x"5F",x"06",x"8C",x"B1",x"91",x"94", -- 0x0420
    x"B8",x"80",x"8C",x"90",x"90",x"90",x"93",x"B6", -- 0x0428
    x"A0",x"B6",x"98",x"96",x"94",x"94",x"93",x"91", -- 0x0430
    x"93",x"93",x"94",x"96",x"B8",x"A0",x"96",x"76", -- 0x0438
    x"74",x"96",x"76",x"74",x"AC",x"B0",x"D1",x"FF", -- 0x0440
    x"1F",x"05",x"5F",x"06",x"80",x"B1",x"B1",x"B1", -- 0x0448
    x"B1",x"AC",x"AC",x"AC",x"AC",x"AA",x"AA",x"AA", -- 0x0450
    x"AA",x"AC",x"AC",x"AC",x"AC",x"8A",x"80",x"8A", -- 0x0458
    x"80",x"AC",x"AC",x"B1",x"FF",x"E7",x"3E",x"01", -- 0x0460
    x"32",x"C8",x"42",x"32",x"C3",x"42",x"F7",x"C3", -- 0x0468
    x"70",x"16",x"DD",x"21",x"B0",x"42",x"DD",x"7E", -- 0x0470
    x"00",x"FE",x"FF",x"28",x"25",x"CD",x"A9",x"14", -- 0x0478
    x"AF",x"C9",x"E7",x"3E",x"00",x"32",x"C3",x"42", -- 0x0480
    x"F7",x"C3",x"6B",x"16",x"3A",x"C8",x"42",x"A7", -- 0x0488
    x"20",x"14",x"E7",x"DD",x"21",x"B0",x"42",x"DD", -- 0x0490
    x"7E",x"00",x"FE",x"FF",x"C8",x"CD",x"A9",x"14", -- 0x0498
    x"AF",x"C9",x"AF",x"32",x"C8",x"42",x"3E",x"FF", -- 0x04A0
    x"C9",x"DD",x"35",x"01",x"C0",x"3A",x"C2",x"42", -- 0x04A8
    x"DD",x"77",x"01",x"DD",x"7E",x"08",x"A7",x"28", -- 0x04B0
    x"16",x"21",x"C4",x"42",x"35",x"7E",x"A7",x"28", -- 0x04B8
    x"0B",x"CD",x"4D",x"02",x"ED",x"5B",x"C5",x"42", -- 0x04C0
    x"19",x"EF",x"18",x"03",x"DD",x"77",x"08",x"DD", -- 0x04C8
    x"CB",x"00",x"46",x"C2",x"E3",x"14",x"DD",x"7E", -- 0x04D0
    x"07",x"D6",x"01",x"FA",x"E3",x"14",x"DD",x"77", -- 0x04D8
    x"07",x"47",x"DF",x"DD",x"35",x"00",x"C0",x"DD", -- 0x04E0
    x"6E",x"02",x"DD",x"66",x"03",x"7E",x"47",x"E6", -- 0x04E8
    x"1F",x"CA",x"94",x"15",x"FE",x"1F",x"C2",x"AE", -- 0x04F0
    x"15",x"23",x"DD",x"75",x"02",x"DD",x"74",x"03", -- 0x04F8
    x"78",x"E6",x"E0",x"0F",x"0F",x"0F",x"0F",x"4F", -- 0x0500
    x"06",x"00",x"21",x"16",x"15",x"09",x"5E",x"23", -- 0x0508
    x"56",x"2A",x"B2",x"42",x"D5",x"C9",x"26",x"15", -- 0x0510
    x"39",x"15",x"49",x"15",x"52",x"15",x"8C",x"15", -- 0x0518
    x"8C",x"15",x"8C",x"15",x"8C",x"15",x"4E",x"CB", -- 0x0520
    x"21",x"CB",x"21",x"06",x"00",x"21",x"E3",x"15", -- 0x0528
    x"09",x"DD",x"75",x"04",x"DD",x"74",x"05",x"18", -- 0x0530
    x"43",x"4E",x"06",x"00",x"21",x"5B",x"16",x"09", -- 0x0538
    x"7E",x"32",x"C2",x"42",x"DD",x"77",x"01",x"18", -- 0x0540
    x"33",x"7E",x"DD",x"77",x"06",x"DD",x"77",x"07", -- 0x0548
    x"18",x"2A",x"7E",x"DD",x"77",x"08",x"DD",x"77", -- 0x0550
    x"09",x"A7",x"28",x"20",x"47",x"E6",x"E0",x"07", -- 0x0558
    x"07",x"07",x"32",x"C4",x"42",x"78",x"16",x"00", -- 0x0560
    x"21",x"00",x"00",x"E6",x"0F",x"87",x"5F",x"78", -- 0x0568
    x"E6",x"10",x"20",x"04",x"ED",x"52",x"18",x"01", -- 0x0570
    x"19",x"22",x"C5",x"42",x"DD",x"6E",x"02",x"DD", -- 0x0578
    x"66",x"03",x"23",x"DD",x"75",x"02",x"DD",x"74", -- 0x0580
    x"03",x"C3",x"E7",x"14",x"06",x"00",x"DF",x"DD", -- 0x0588
    x"36",x"00",x"FF",x"C9",x"CD",x"9C",x"15",x"06", -- 0x0590
    x"00",x"DF",x"18",x"39",x"78",x"E6",x"E0",x"07", -- 0x0598
    x"07",x"07",x"47",x"3E",x"01",x"10",x"04",x"DD", -- 0x05A0
    x"77",x"00",x"C9",x"07",x"18",x"F7",x"C5",x"CD", -- 0x05A8
    x"9C",x"15",x"C1",x"78",x"E6",x"1F",x"3D",x"07", -- 0x05B0
    x"4F",x"06",x"00",x"DD",x"6E",x"04",x"DD",x"66", -- 0x05B8
    x"05",x"09",x"5E",x"23",x"56",x"EB",x"EF",x"DD", -- 0x05C0
    x"7E",x"09",x"DD",x"77",x"08",x"DD",x"46",x"06", -- 0x05C8
    x"78",x"DD",x"77",x"07",x"DF",x"DD",x"6E",x"02", -- 0x05D0
    x"DD",x"66",x"03",x"23",x"DD",x"75",x"02",x"DD", -- 0x05D8
    x"74",x"03",x"C9",x"6B",x"08",x"F2",x"07",x"80", -- 0x05E0
    x"07",x"14",x"07",x"AE",x"06",x"4E",x"06",x"F3", -- 0x05E8
    x"05",x"9E",x"05",x"4E",x"05",x"01",x"05",x"B9", -- 0x05F0
    x"04",x"76",x"04",x"36",x"04",x"F9",x"03",x"C0", -- 0x05F8
    x"03",x"8A",x"03",x"57",x"03",x"27",x"03",x"FA", -- 0x0600
    x"02",x"CF",x"02",x"A7",x"02",x"81",x"02",x"5D", -- 0x0608
    x"02",x"3B",x"02",x"1B",x"02",x"FD",x"01",x"E0", -- 0x0610
    x"01",x"C5",x"01",x"AC",x"01",x"94",x"01",x"7D", -- 0x0618
    x"01",x"68",x"01",x"53",x"01",x"40",x"01",x"2E", -- 0x0620
    x"01",x"1D",x"01",x"0D",x"01",x"FE",x"00",x"F0", -- 0x0628
    x"00",x"E3",x"00",x"D6",x"00",x"CA",x"00",x"BE", -- 0x0630
    x"00",x"B4",x"00",x"AA",x"00",x"A0",x"00",x"97", -- 0x0638
    x"00",x"8F",x"00",x"87",x"00",x"7F",x"00",x"78", -- 0x0640
    x"00",x"71",x"00",x"6B",x"00",x"65",x"00",x"5F", -- 0x0648
    x"00",x"5A",x"00",x"55",x"00",x"50",x"00",x"4C", -- 0x0650
    x"00",x"47",x"00",x"11",x"0F",x"0D",x"0B",x"0A", -- 0x0658
    x"09",x"08",x"07",x"03",x"05",x"14",x"13",x"11", -- 0x0660
    x"10",x"0F",x"0E",x"3A",x"C8",x"42",x"A7",x"C0", -- 0x0668
    x"21",x"94",x"16",x"11",x"B0",x"42",x"01",x"0A", -- 0x0670
    x"00",x"ED",x"B0",x"3A",x"C3",x"42",x"87",x"4F", -- 0x0678
    x"87",x"81",x"4F",x"21",x"9E",x"16",x"09",x"11", -- 0x0680
    x"B2",x"42",x"7E",x"12",x"CD",x"91",x"16",x"7E", -- 0x0688
    x"12",x"23",x"13",x"C9",x"01",x"01",x"00",x"00", -- 0x0690
    x"00",x"00",x"00",x"00",x"00",x"00",x"AA",x"16", -- 0x0698
    x"CD",x"16",x"CD",x"16",x"B8",x"16",x"CD",x"16", -- 0x06A0
    x"CD",x"16",x"1F",x"0F",x"3F",x"09",x"5F",x"09", -- 0x06A8
    x"7F",x"00",x"6D",x"71",x"74",x"79",x"D6",x"FF", -- 0x06B0
    x"1F",x"02",x"3F",x"07",x"5F",x"09",x"7F",x"00", -- 0x06B8
    x"94",x"8D",x"88",x"94",x"8D",x"88",x"94",x"8D", -- 0x06C0
    x"88",x"94",x"8D",x"C8",x"FF",x"FF",x"FF",x"FF", -- 0x06C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x07F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
