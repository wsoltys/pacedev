`timescale 1ns / 1ps
module COCO3VIDEO(
PIX_CLK,
RESET_N,
RED1,
GREEN1,
BLUE1,
RED0,
GREEN0,
BLUE0,
HSYNC,
SYNC_FLAG,
VSYNC,
READMEM,
RAM_ADDRESS,
RAM_DATA,
VBANK,
COCO,
V,
BP,
VERT,
VID_CONT,
CSS,
LPF,
VERT_FIN_SCRL,
LPR,
HRES,
CRES,
HVEN,
HOR_OFFSET,
SCRN_START_MSB,
SCRN_START_LSB,
BDR_PAL,
PALETTE0,
PALETTE1,
PALETTE2,
PALETTE3,
PALETTE4,
PALETTE5,
PALETTE6,
PALETTE7,
PALETTE8,
PALETTE9,
PALETTEA,
PALETTEB,
PALETTEC,
PALETTED,
PALETTEE,
PALETTEF,
BLINK
);

input					PIX_CLK;
input					RESET_N;
output				RED1;
output				GREEN1;
output				BLUE1;
output				RED0;
output				GREEN0;
output				BLUE0;
reg					RED1;
reg					GREEN1;
reg					BLUE1;
reg					RED0;
reg					GREEN0;
reg					BLUE0;
output				HSYNC;
reg					HSYNC;
output				SYNC_FLAG;
reg					SYNC_FLAG;
output				VSYNC;
reg					VSYNC;
output				READMEM;
reg					READMEM;
output	[17:0]	RAM_ADDRESS;
input		[31:0]	RAM_DATA;
input					VBANK;
input					COCO;
input		[2:0]		V;
input					BP;
input		[6:0]		VERT;
input		[3:0]		VID_CONT;
input					CSS;
input		[1:0]		LPF;
input		[2:0]		LPR;
input		[3:0]		VERT_FIN_SCRL;
input		[2:0]		HRES;
input		[1:0]		CRES;
input					HVEN;
input		[6:0]		HOR_OFFSET;
input		[7:0]		SCRN_START_MSB;
input		[7:0]		SCRN_START_LSB;
input		[5:0]		BDR_PAL;
input		[5:0]		PALETTE0;
input		[5:0]		PALETTE1;
input		[5:0]		PALETTE2;
input		[5:0]		PALETTE3;
input		[5:0]		PALETTE4;
input		[5:0]		PALETTE5;
input		[5:0]		PALETTE6;
input		[5:0]		PALETTE7;
input		[5:0]		PALETTE8;
input		[5:0]		PALETTE9;
input		[5:0]		PALETTEA;
input		[5:0]		PALETTEB;
input		[5:0]		PALETTEC;
input		[5:0]		PALETTED;
input		[5:0]		PALETTEE;
input		[5:0]		PALETTEF;
input					BLINK;

reg		[9:0]		LINE;
reg		[4:0]		VLPR;
reg		[7:0]		VADD;
reg		[9:0]		PIXEL_COUNT;
reg		[7:0]		CHAR_LATCH;
reg		[7:0]		CHAR_LATCH3;
reg		[7:0]		ATRIB_LATCH;
reg		[7:0]		ATRIB_LATCH3;
wire		[3:0]		PIXEL_ORDER;
reg					HBLANKING;
reg					VBLANKING;
wire					READROM1;
wire					READROM2;
reg		[7:0]		CHARACTER;
wire		[7:0]		CHARACTER1;
reg		[7:0]		CHARACTER2;
reg		[7:0]		CHARACTER3;
wire		[7:0]		CHARACTER4;
reg					ROW;
wire					MODE_256;
wire					COCO_GR;
wire					BLINK;

wire		[10:0]	ROM_ADDRESS;
wire		[7:0]		ROM_DATA1;
wire		[2:0]		LINES_ROW;
reg					SIX;
wire					RED1X;
wire					GREEN1X;
wire					BLUE1X;
wire					RED0X;
wire					GREEN0X;
wire					BLUE0X;
wire		[5:0]		PIXEL0;
wire		[5:0]		PIXEL1;
wire		[5:0]		PIXEL2;
wire		[5:0]		PIXEL3;
wire		[5:0]		PIXEL4;
wire		[5:0]		PIXEL5;
wire		[5:0]		PIXEL6;
wire		[5:0]		PIXEL7;
wire		[5:0]		PIXEL8;
wire		[5:0]		PIXEL9;
wire		[5:0]		PIXELA;
wire		[5:0]		PIXELB;
wire		[5:0]		PIXELC;
wire		[5:0]		PIXELD;
wire		[5:0]		PIXELE;
wire		[5:0]		PIXELF;
reg		[15:0]	RED1S;
reg		[15:0]	RED0S;
reg		[15:0]	GREEN1S;
reg		[15:0]	GREEN0S;
reg		[15:0]	BLUE1S;
reg		[15:0]	BLUE0S;
reg		[18:0]	ROW_ADD;
wire		[18:0]	START_ADD;
reg					VBORDER;
reg					HBORDER;
wire		[5:0]		BORDER;

// Character generator
`include "COCO3GEN.v"

/*****************************************************************************
* Generate master pixel clock
******************************************************************************/
//always @(posedge CLK)
//begin
//		PIX_CLK <= ~PIX_CLK;
//end
/*****************************************************************************
* Read RAM
******************************************************************************/
assign RAM_ADDRESS =
// CoCo1 low res graphics (64 pixels / 2 bytes)
({COCO,V[0]} == 2'b11)						?	ROW_ADD[18:1] + PIXEL_COUNT[9:6]:
//	HR Text
({COCO,BP,HRES[2],CRES[0]}==4'b0000)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:5]:	//32 / 40
({COCO,BP,HRES[2],CRES[0]}==4'b0001)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:4]:	//64 / 80
({COCO,BP,HRES[2],CRES[0]}==4'b0010)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:4]:	//64 / 80
({COCO,BP,HRES[2],CRES[0]}==4'b0011)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:3]:	//128 /160
//	HR Graphics
							({COCO,BP,HRES}==5'b01000)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:6]:	//16
							({COCO,BP,HRES}==5'b01001)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:6]:	//20
							({COCO,BP,HRES}==5'b01010)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:5]:	//32
							({COCO,BP,HRES}==5'b01011)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:5]:	//40
							({COCO,BP,HRES}==5'b01100)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:4]:	//64
							({COCO,BP,HRES}==5'b01101)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:4]:	//80
							({COCO,BP,HRES}==5'b01110)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:3]:	//128
							({COCO,BP,HRES}==5'b01111)	?	ROW_ADD[18:1] + PIXEL_COUNT[9:3]:	//160
// CoCo1 Text
																	ROW_ADD[18:1] + PIXEL_COUNT[9:5];	//32

//HVEN,
//HOR_OFFSET,
//input		[7:0]		SCRN_START_MSB;
//input		[7:0]		SCRN_START_LSB;
assign START_ADD =
// CoCo1 low res graphics (64 pixels / 2 bytes)
({COCO,V[0]} == 2'b11)										?	ROW_ADD + 9'd16:
// HR Text
({HVEN,COCO} == 2'b10)										?  ROW_ADD + 9'd256:
({HVEN,COCO,BP,HRES[2],CRES[0],HRES[0]}==6'b000000)?	ROW_ADD + 9'd32:
({HVEN,COCO,BP,HRES[2],CRES[0],HRES[0]}==6'b000001)?	ROW_ADD + 9'd40:
({HVEN,COCO,BP,HRES[2],CRES[0],HRES[0]}==6'b000010)?	ROW_ADD + 9'd64:
({HVEN,COCO,BP,HRES[2],CRES[0],HRES[0]}==6'b000011)?	ROW_ADD + 9'd80:
({HVEN,COCO,BP,HRES[2],CRES[0],HRES[0]}==6'b000100)?	ROW_ADD + 9'd64:
({HVEN,COCO,BP,HRES[2],CRES[0],HRES[0]}==6'b000101)?	ROW_ADD + 9'd80:
({HVEN,COCO,BP,HRES[2],CRES[0],HRES[0]}==6'b000110)?	ROW_ADD + 9'd128:
({HVEN,COCO,BP,HRES[2],CRES[0],HRES[0]}==6'b000111)?	ROW_ADD + 9'd160:
//	HR Graphics
						({HVEN,COCO,BP,HRES}==6'b001000)	?	ROW_ADD + 9'd16:
						({HVEN,COCO,BP,HRES}==6'b001001)	?	ROW_ADD + 9'd20:
						({HVEN,COCO,BP,HRES}==6'b001010)	?	ROW_ADD + 9'd32:
						({HVEN,COCO,BP,HRES}==6'b001011)	?	ROW_ADD + 9'd40:
						({HVEN,COCO,BP,HRES}==6'b001100)	?	ROW_ADD + 9'd64:
						({HVEN,COCO,BP,HRES}==6'b001101)	?	ROW_ADD + 9'd80:
						({HVEN,COCO,BP,HRES}==6'b001110)	?	ROW_ADD + 9'd128:
						({HVEN,COCO,BP,HRES}==6'b001111)	?	ROW_ADD + 9'd160:
// CoCo1 Text
																		ROW_ADD + 9'd32;

//assign READMEM =	(PIXEL_COUNT[2:0] == 3'b000)									?	1'b1:
//						(PIXEL_COUNT[2:0] == 3'b001)									?	1'b1:
//			 																						1'b0;

/*****************************************************************************
* Read Character ROM
******************************************************************************/
//VID_CONT[0] will change to lower case mode in coco1=1 mode
//VID_CONT[1] will invert forground and background in coco1=1 mode
assign ROM_ADDRESS =	({COCO,PIXEL_COUNT[2],VID_CONT[0]} == 3'b100)							?	{~CHAR_LATCH[5], CHAR_LATCH[5:0], VLPR[4:1]}:	// COCO1 Text 1 w/o LC
							({COCO,PIXEL_COUNT[2],VID_CONT[0]} == 3'b110)							?	{~ATRIB_LATCH[5], ATRIB_LATCH[5:0], VLPR[4:1]}:	// COCO1 Text 2 w/o LC
							({COCO,PIXEL_COUNT[2],VID_CONT[0],CHAR_LATCH[6]} == 4'b1011)		?	{~CHAR_LATCH[5], CHAR_LATCH[5:0], VLPR[4:1]}:	// COCO1 Text 1 w/o LC
							({COCO,PIXEL_COUNT[2],VID_CONT[0],ATRIB_LATCH[6]} == 4'b1111)		?	{~ATRIB_LATCH[5], ATRIB_LATCH[5:0], VLPR[4:1]}:	// COCO1 Text 2 w/o LC
							({COCO,PIXEL_COUNT[2],VID_CONT[0],CHAR_LATCH[6:5]} == 5'b10101)	?	{~CHAR_LATCH[5], CHAR_LATCH[5:0], VLPR[4:1]}:	// COCO1 Text 1 w/o LC
							({COCO,PIXEL_COUNT[2],VID_CONT[0],ATRIB_LATCH[6:5]} == 5'b11101)	?	{~ATRIB_LATCH[5], ATRIB_LATCH[5:0], VLPR[4:1]}:	// COCO1 Text 2 w/o LC
							({COCO,PIXEL_COUNT[2],VID_CONT[0],CHAR_LATCH[6:5]} == 5'b10100)	?	{2'b11, CHAR_LATCH[4:0], VLPR[4:1]}:	// COCO1 Text 1 with LC
							({COCO,PIXEL_COUNT[2],VID_CONT[0],ATRIB_LATCH[6:5]} == 5'b11100)	?	{2'b11, ATRIB_LATCH[4:0], VLPR[4:1]}:	// COCO1 Text 2 with LC
							({COCO,PIXEL_COUNT[2]} == 2'b00)												?	{CHAR_LATCH[6:0], VLPR[4:1]}:		// COCO3 Text 1
																														{ATRIB_LATCH[6:0], VLPR[4:1]};		// COCO3 Text 2

assign READROM1 =	(PIXEL_COUNT[2:0] == 3'b010)			?	1'b1:
																			1'b0;

always @(negedge READROM1)
begin
	if({COCO,BP,CRES[0],ATRIB_LATCH[6],ROW,SIX} == 6'b001111)
		CHARACTER <=	8'hFF;
	else
		CHARACTER <=	ROM_DATA1;

		CHARACTER3 <=	CHARACTER1;
end

assign CHARACTER1 =	({COCO,BP,CRES[0],ATRIB_LATCH[7],BLINK} == 5'b00111)	?	8'h00:			// Hires Text blink
							({COCO, VID_CONT[1:0], CHAR_LATCH[6:5]} == 5'b10000)	?	~CHARACTER:		// Lowres  0-31 Normal UC only (Inverse)
							({COCO, VID_CONT[1:0], CHAR_LATCH[6:5]} == 5'b10001)	?	~CHARACTER:		// Lowres 32-64 Normal UC only (Inverse)
							({COCO, VID_CONT[1:0], CHAR_LATCH[6:5]} == 5'b10101)	?	~CHARACTER:		// Lowres 32-64 LC but UC part (Inverse)
							({COCO, VID_CONT[1:0], CHAR_LATCH[6:5]} == 5'b11010)	?	~CHARACTER:		// Lowres 64-95 Inverse
							({COCO, VID_CONT[1:0], CHAR_LATCH[6:5]} == 5'b11011)	?	~CHARACTER:		// Lowres 96-128 Inverse
							({COCO, VID_CONT[1:0], CHAR_LATCH[6:5]} == 5'b11100)	?	~CHARACTER:		// Lowres  0-31 Inverse
							({COCO, VID_CONT[1:0], CHAR_LATCH[6:5]} == 5'b11110)	?	~CHARACTER:		// Lowres 64-95 Inverse
							({COCO, VID_CONT[1:0], CHAR_LATCH[6:5]} == 5'b11111)	?	~CHARACTER:		// Lowres 96-128 Inverse
																										 CHARACTER;		// Normal Video

assign READROM2 =	(PIXEL_COUNT[2:0] == 3'b110)			?	1'b1:
																			1'b0;

assign CHARACTER4 =	({COCO, VID_CONT[1:0], ATRIB_LATCH[6:5]} == 5'b10000)	?	~CHARACTER2:		// Lowres  0-31 Normal UC only (Inverse)
							({COCO, VID_CONT[1:0], ATRIB_LATCH[6:5]} == 5'b10001)	?	~CHARACTER2:		// Lowres 32-64 Normal UC only (Inverse)
							({COCO, VID_CONT[1:0], ATRIB_LATCH[6:5]} == 5'b10101)	?	~CHARACTER2:		// Lowres 32-64 LC but UC part (Inverse)
							({COCO, VID_CONT[1:0], ATRIB_LATCH[6:5]} == 5'b11010)	?	~CHARACTER2:		// Lowres 64-95 Inverse
							({COCO, VID_CONT[1:0], ATRIB_LATCH[6:5]} == 5'b11011)	?	~CHARACTER2:		// Lowres 96-128 Inverse
							({COCO, VID_CONT[1:0], ATRIB_LATCH[6:5]} == 5'b11100)	?	~CHARACTER2:		// Lowres  0-31 Inverse
							({COCO, VID_CONT[1:0], ATRIB_LATCH[6:5]} == 5'b11110)	?	~CHARACTER2:		// Lowres 64-95 Inverse
							({COCO, VID_CONT[1:0], ATRIB_LATCH[6:5]} == 5'b11111)	?	~CHARACTER2:		// Lowres 96-128 Inverse
																										 CHARACTER2;		// Normal Video

always @(negedge READROM2)
begin
	CHARACTER2 <=	ROM_DATA1;
end

assign	COCO_GR	=	(V == 3'b000)		?	1'b0:
//							(COCO == 1'b0)		?	1'b0:
														1'b1;
assign PIXEL0 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,CHAR_LATCH[7],CHARACTER1[0]} == 6'b100001)			?	PALETTEC:
			({COCO,V,CHAR_LATCH[7],CHARACTER1[0]} == 6'b100000)			?	PALETTED:
//			({COCO,V,CHAR_LATCH[7,6],CHARACTER1[0]} == 7'b1000010)			?	PALETTED:
//			({COCO,V,CHAR_LATCH[7,6],CHARACTER1[0]} == 7'b1000011)			?	PALETTEC:
// HR Text 80 (2 bytes is 1-8 pixel character)
// HR Text 40 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[5:3]}==7'b0011000)	?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[5:3]}==7'b0011001)	?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[5:3]}==7'b0011010)	?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[5:3]}==7'b0011011)	?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[5:3]}==7'b0011100)	?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[5:3]}==7'b0011101)	?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[5:3]}==7'b0011110)	?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[5:3]}==7'b0011111)	?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[2:0]}==7'b0010000)	?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[2:0]}==7'b0010001)	?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[2:0]}==7'b0010010)	?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[2:0]}==7'b0010011)	?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[2:0]}==7'b0010100)	?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[2:0]}==7'b0010101)	?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[2:0]}==7'b0010110)	?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER1[0],ATRIB_LATCH[2:0]}==7'b0010111)	?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER1[0]}==4'b0001)							?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[0]}==4'b0000)							?	PALETTED:
//SG4 (2 bytes is 2-8 (really 2) pixels)
			({COCO,V,CHAR_LATCH[7],SIX,  CHAR_LATCH[0]} == 7'b1000110)				?	PALETTE8:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[0]} == 10'b1000100011)			?	PALETTE0:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[0]} == 10'b1000100111)			?	PALETTE1:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[0]} == 10'b1000101011)			?	PALETTE2:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[0]} == 10'b1000101111)			?	PALETTE3:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[0]} == 10'b1000110011)			?	PALETTE4:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[0]} == 10'b1000110111)			?	PALETTE5:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[0]} == 10'b1000111011)			?	PALETTE6:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[0]} == 10'b1000111111)			?	PALETTE7:
			({COCO,V,CHAR_LATCH[7],SIX,  CHAR_LATCH[2]} == 7'b1000100)				?	PALETTE8:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[2]} == 10'b1000100001)			?	PALETTE0:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[2]} == 10'b1000100101)			?	PALETTE1:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[2]} == 10'b1000101001)			?	PALETTE2:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[2]} == 10'b1000101101)			?	PALETTE3:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[2]} == 10'b1000110001)			?	PALETTE4:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[2]} == 10'b1000110101)			?	PALETTE5:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[2]} == 10'b1000111001)			?	PALETTE6:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[2]} == 10'b1000111101)			?	PALETTE7:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[0]} == 5'b11100)		?	PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[0]} == 5'b11101)		?	PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[0]} == 5'b11110)		?	PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[0]} == 5'b11111)		?	PALETTEB:
// 4 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1:0]} == 6'b110000)	?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1:0]} == 6'b110001)	?	PALETTE1:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1:0]} == 6'b110010)	?	PALETTE2:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1:0]} == 6'b110011)	?	PALETTE3:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1:0]} == 6'b110100)	?	PALETTE4:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1:0]} == 6'b110101)	?	PALETTE5:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1:0]} == 6'b110110)	?	PALETTE6:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1:0]} == 6'b110111)	?	PALETTE7:
// Hires GR
// 2 color
			({COCO,BP,CRES,CHAR_LATCH[0]} == 5'b01000)							?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[0]} == 5'b01001)							?	PALETTE1:
// 4 Color
			({COCO,BP,CRES,CHAR_LATCH[1:0]} == 6'b010100)						?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[1:0]} == 6'b010101)						?	PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH[1:0]} == 6'b010110)						?	PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH[1:0]} == 6'b010111)						?	PALETTE3:
// 16 color
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01100000)						?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01100001)						?	PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01100010)						?	PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01100011)						?	PALETTE3:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01100100)						?	PALETTE4:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01100101)						?	PALETTE5:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01100110)						?	PALETTE6:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01100111)						?	PALETTE7:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01101000)						?	PALETTE8:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01101001)						?	PALETTE9:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01101010)						?	PALETTEA:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01101011)						?	PALETTEB:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01101100)						?	PALETTEC:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01101101)						?	PALETTED:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01101110)						?	PALETTEE:
			({COCO,BP,CRES,CHAR_LATCH[3:0]} == 8'b01101111)						?	PALETTEF:
																									PALETTE0;

assign PIXEL1 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,CHAR_LATCH[7],CHARACTER1[1]} == 6'b100001)			?	PALETTEC:
			({COCO,V,CHAR_LATCH[7],CHARACTER1[1]} == 6'b100000)			?	PALETTED:
// HR Text 80 (2 bytes is 1-8 pixel character)
// HR Text 40 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[5:3]}==7'b0011000)	?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[5:3]}==7'b0011001)	?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[5:3]}==7'b0011010)	?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[5:3]}==7'b0011011)	?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[5:3]}==7'b0011100)	?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[5:3]}==7'b0011101)	?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[5:3]}==7'b0011110)	?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[5:3]}==7'b0011111)	?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[2:0]}==7'b0010000)	?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[2:0]}==7'b0010001)	?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[2:0]}==7'b0010010)	?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[2:0]}==7'b0010011)	?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[2:0]}==7'b0010100)	?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[2:0]}==7'b0010101)	?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[2:0]}==7'b0010110)	?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER1[1],ATRIB_LATCH[2:0]}==7'b0010111)	?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER1[1]}==4'b0001)							?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[1]}==4'b0000)							?	PALETTED:
//SG4 (2 bytes is 2-8 (really 2) pixels)
			({COCO,V,CHAR_LATCH[7],SIX,  CHAR_LATCH[1]} == 7'b1000110)				?	PALETTE8:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[1]} == 10'b1000100011)			?	PALETTE0:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[1]} == 10'b1000100111)			?	PALETTE1:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[1]} == 10'b1000101011)			?	PALETTE2:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[1]} == 10'b1000101111)			?	PALETTE3:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[1]} == 10'b1000110011)			?	PALETTE4:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[1]} == 10'b1000110111)			?	PALETTE5:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[1]} == 10'b1000111011)			?	PALETTE6:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[1]} == 10'b1000111111)			?	PALETTE7:
			({COCO,V,CHAR_LATCH[7],SIX,  CHAR_LATCH[3]} == 7'b1000100)				?	PALETTE8:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[3]} == 10'b1000100001)			?	PALETTE0:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[3]} == 10'b1000100101)			?	PALETTE1:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[3]} == 10'b1000101001)			?	PALETTE2:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[3]} == 10'b1000101101)			?	PALETTE3:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[3]} == 10'b1000110001)			?	PALETTE4:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[3]} == 10'b1000110101)			?	PALETTE5:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[3]} == 10'b1000111001)			?	PALETTE6:
			({COCO,V,CHAR_LATCH[7:4],SIX,CHAR_LATCH[3]} == 10'b1000111101)			?	PALETTE7:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1]} == 5'b11100)		?	PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1]} == 5'b11101)		?	PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1]} == 5'b11110)		?	PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[1]} == 5'b11111)		?	PALETTEB:
// 4 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3:2]} == 6'b110000)	?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3:2]} == 6'b110001)	?	PALETTE1:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3:2]} == 6'b110010)	?	PALETTE2:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3:2]} == 6'b110011)	?	PALETTE3:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3:2]} == 6'b110100)	?	PALETTE4:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3:2]} == 6'b110101)	?	PALETTE5:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3:2]} == 6'b110110)	?	PALETTE6:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3:2]} == 6'b110111)	?	PALETTE7:
// Hires GR
// 2 color
			({COCO,BP,CRES,CHAR_LATCH[1]} == 5'b01000)							?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[1]} == 5'b01001)							?	PALETTE1:
// 4 Color
			({COCO,BP,CRES,CHAR_LATCH[3:2]} == 6'b010100)						?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[3:2]} == 6'b010101)						?	PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH[3:2]} == 6'b010110)						?	PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH[3:2]} == 6'b010111)						?	PALETTE3:
// 16 color
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01100000)						?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01100001)						?	PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01100010)						?	PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01100011)						?	PALETTE3:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01100100)						?	PALETTE4:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01100101)						?	PALETTE5:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01100110)						?	PALETTE6:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01100111)						?	PALETTE7:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01101000)						?	PALETTE8:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01101001)						?	PALETTE9:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01101010)						?	PALETTEA:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01101011)						?	PALETTEB:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01101100)						?	PALETTEC:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01101101)						?	PALETTED:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01101110)						?	PALETTEE:
			({COCO,BP,CRES,CHAR_LATCH[7:4]} == 8'b01101111)						?	PALETTEF:
																									PALETTE0;

assign PIXEL2 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,CHAR_LATCH[7],CHARACTER1[2],PIXEL_COUNT[4]} == 7'b1000010)			?	PALETTEC:
			({COCO,V,CHAR_LATCH[7],CHARACTER1[2],PIXEL_COUNT[4]} == 7'b1000000)			?	PALETTED:
// HR Text 80 (2 bytes is 1-8 pixel character)
// HR Text 40 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[5:3]}==7'b0011000)	?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[5:3]}==7'b0011001)	?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[5:3]}==7'b0011010)	?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[5:3]}==7'b0011011)	?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[5:3]}==7'b0011100)	?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[5:3]}==7'b0011101)	?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[5:3]}==7'b0011110)	?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[5:3]}==7'b0011111)	?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[2:0]}==7'b0010000)	?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[2:0]}==7'b0010001)	?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[2:0]}==7'b0010010)	?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[2:0]}==7'b0010011)	?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[2:0]}==7'b0010100)	?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[2:0]}==7'b0010101)	?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[2:0]}==7'b0010110)	?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER1[2],ATRIB_LATCH[2:0]}==7'b0010111)	?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER1[2]}==4'b0001)							?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[2]}==4'b0000)							?	PALETTED:
//SG4 (2 bytes is 2-8 (really 2) pixels)
			({COCO,V,ATRIB_LATCH[7],SIX,  ATRIB_LATCH[0]} == 7'b1000110)			?	PALETTE8:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[0]} == 10'b1000100011)		?	PALETTE0:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[0]} == 10'b1000100111)		?	PALETTE1:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[0]} == 10'b1000101011)		?	PALETTE2:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[0]} == 10'b1000101111)		?	PALETTE3:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[0]} == 10'b1000110011)		?	PALETTE4:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[0]} == 10'b1000110111)		?	PALETTE5:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[0]} == 10'b1000111011)		?	PALETTE6:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[0]} == 10'b1000111111)		?	PALETTE7:
			({COCO,V,ATRIB_LATCH[7],SIX,  ATRIB_LATCH[2]} == 7'b1000100)			?	PALETTE8:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[2]} == 10'b1000100001)		?	PALETTE0:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[2]} == 10'b1000100101)		?	PALETTE1:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[2]} == 10'b1000101001)		?	PALETTE2:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[2]} == 10'b1000101101)		?	PALETTE3:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[2]} == 10'b1000110001)		?	PALETTE4:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[2]} == 10'b1000110101)		?	PALETTE5:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[2]} == 10'b1000111001)		?	PALETTE6:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[2]} == 10'b1000111101)		?	PALETTE7:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[2]} == 5'b11100)		?	PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[2]} == 5'b11101)		?	PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[2]} == 5'b11110)		?	PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[2]} == 5'b11111)		?	PALETTEB:
// 4 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5:4]} == 6'b110000)	?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5:4]} == 6'b110001)	?	PALETTE1:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5:4]} == 6'b110010)	?	PALETTE2:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5:4]} == 6'b110011)	?	PALETTE3:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5:4]} == 6'b110100)	?	PALETTE4:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5:4]} == 6'b110101)	?	PALETTE5:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5:4]} == 6'b110110)	?	PALETTE6:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5:4]} == 6'b110111)	?	PALETTE7:
// Hires GR
// 2 color
			({COCO,BP,CRES,CHAR_LATCH[2]} == 5'b01000)							?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[2]} == 5'b01001)							?	PALETTE1:
// 4 Color
			({COCO,BP,CRES,CHAR_LATCH[5:4]} == 6'b010100)						?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[5:4]} == 6'b010101)						?	PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH[5:4]} == 6'b010110)						?	PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH[5:4]} == 6'b010111)						?	PALETTE3:
// 16 color
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01100000)					?	PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01100001)					?	PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01100010)					?	PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01100011)					?	PALETTE3:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01100100)					?	PALETTE4:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01100101)					?	PALETTE5:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01100110)					?	PALETTE6:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01100111)					?	PALETTE7:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01101000)					?	PALETTE8:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01101001)					?	PALETTE9:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01101010)					?	PALETTEA:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01101011)					?	PALETTEB:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01101100)					?	PALETTEC:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01101101)					?	PALETTED:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01101110)					?	PALETTEE:
			({COCO,BP,CRES,ATRIB_LATCH[3:0]} == 8'b01101111)					?	PALETTEF:
																									PALETTE0;

assign PIXEL3 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,CHAR_LATCH[7],CHARACTER1[3],PIXEL_COUNT[4]} == 7'b1000010)			?	PALETTEC:
			({COCO,V,CHAR_LATCH[7],CHARACTER1[3],PIXEL_COUNT[4]} == 7'b1000000)			?	PALETTED:
// HR Text 80 (2 bytes is 1-8 pixel character)
// HR Text 40 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[5:3]}==7'b0011000)	?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[5:3]}==7'b0011001)	?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[5:3]}==7'b0011010)	?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[5:3]}==7'b0011011)	?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[5:3]}==7'b0011100)	?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[5:3]}==7'b0011101)	?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[5:3]}==7'b0011110)	?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[5:3]}==7'b0011111)	?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[2:0]}==7'b0010000)	?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[2:0]}==7'b0010001)	?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[2:0]}==7'b0010010)	?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[2:0]}==7'b0010011)	?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[2:0]}==7'b0010100)	?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[2:0]}==7'b0010101)	?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[2:0]}==7'b0010110)	?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER1[3],ATRIB_LATCH[2:0]}==7'b0010111)	?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER1[3]}==4'b0001)							?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[3]}==4'b0000)							?	PALETTED:
//SG4 (2 bytes is 2-8 (really 2) pixels)
			({COCO,V,ATRIB_LATCH[7],SIX,  ATRIB_LATCH[1]} == 7'b1000110)			?	PALETTE8:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[1]} == 10'b1000100011)		?	PALETTE0:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[1]} == 10'b1000100111)		?	PALETTE1:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[1]} == 10'b1000101011)		?	PALETTE2:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[1]} == 10'b1000101111)		?	PALETTE3:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[1]} == 10'b1000110011)		?	PALETTE4:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[1]} == 10'b1000110111)		?	PALETTE5:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[1]} == 10'b1000111011)		?	PALETTE6:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[1]} == 10'b1000111111)		?	PALETTE7:
			({COCO,V,ATRIB_LATCH[7],SIX,  ATRIB_LATCH[3]} == 7'b1000100)			?	PALETTE8:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[3]} == 10'b1000100001)		?	PALETTE0:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[3]} == 10'b1000100101)		?	PALETTE1:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[3]} == 10'b1000101001)		?	PALETTE2:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[3]} == 10'b1000101101)		?	PALETTE3:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[3]} == 10'b1000110001)		?	PALETTE4:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[3]} == 10'b1000110101)		?	PALETTE5:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[3]} == 10'b1000111001)		?	PALETTE6:
			({COCO,V,ATRIB_LATCH[7:4],SIX,ATRIB_LATCH[3]} == 10'b1000111101)		?	PALETTE7:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3]} == 5'b11100)		?	PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3]} == 5'b11101)		?	PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3]} == 5'b11110)		?	PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[3]} == 5'b11111)		?	PALETTEB:
// 4 COLOR
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7:6]} == 6'b110000)	?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7:6]} == 6'b110001)	?	PALETTE1:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7:6]} == 6'b110010)	?	PALETTE2:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7:6]} == 6'b110011)	?	PALETTE3:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7:6]} == 6'b110100)	?	PALETTE4:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7:6]} == 6'b110101)	?	PALETTE5:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7:6]} == 6'b110110)	?	PALETTE6:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7:6]} == 6'b110111)	?	PALETTE7:
// Hires GR
// 2 color
			({COCO,BP,CRES,CHAR_LATCH[3]} == 5'b01000)							?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[3]} == 5'b01001)							?	PALETTE1:
// 4 Color
			({COCO,BP,CRES,CHAR_LATCH[7:6]} == 6'b010100)						?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[7:6]} == 6'b010101)						?	PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH[7:6]} == 6'b010110)						?	PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH[7:6]} == 6'b010111)						?	PALETTE3:
// 16 color
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01100000)					?	PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01100001)					?	PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01100010)					?	PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01100011)					?	PALETTE3:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01100100)					?	PALETTE4:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01100101)					?	PALETTE5:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01100110)					?	PALETTE6:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01100111)					?	PALETTE7:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01101000)					?	PALETTE8:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01101001)					?	PALETTE9:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01101010)					?	PALETTEA:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01101011)					?	PALETTEB:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01101100)					?	PALETTEC:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01101101)					?	PALETTED:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01101110)					?	PALETTEE:
			({COCO,BP,CRES,ATRIB_LATCH[7:4]} == 8'b01101111)					?	PALETTEF:
																									PALETTE0;

assign PIXEL4 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,CHAR_LATCH[7],CHARACTER1[4]} == 6'b100001)			?	PALETTEC:
			({COCO,V,CHAR_LATCH[7],CHARACTER1[4]} == 6'b100000)			?	PALETTED:
// HR Text 80 (2 bytes is 1-8 pixel character)
// HR Text 40 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[5:3]}==7'b0011000)	?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[5:3]}==7'b0011001)	?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[5:3]}==7'b0011010)	?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[5:3]}==7'b0011011)	?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[5:3]}==7'b0011100)	?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[5:3]}==7'b0011101)	?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[5:3]}==7'b0011110)	?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[5:3]}==7'b0011111)	?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[2:0]}==7'b0010000)	?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[2:0]}==7'b0010001)	?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[2:0]}==7'b0010010)	?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[2:0]}==7'b0010011)	?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[2:0]}==7'b0010100)	?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[2:0]}==7'b0010101)	?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[2:0]}==7'b0010110)	?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER1[4],ATRIB_LATCH[2:0]}==7'b0010111)	?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER1[4]}==4'b0001)							?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[4]}==4'b0000)							?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[4]} == 5'b11100)		?	PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[4]} == 5'b11101)		?	PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[4]} == 5'b11110)		?	PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[4]} == 5'b11111)		?	PALETTEB:
// 4 COLOR
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1:0]} == 6'b110000)	?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1:0]} == 6'b110001)	?	PALETTE1:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1:0]} == 6'b110010)	?	PALETTE2:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1:0]} == 6'b110011)	?	PALETTE3:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1:0]} == 6'b110100)	?	PALETTE4:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1:0]} == 6'b110101)	?	PALETTE5:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1:0]} == 6'b110110)	?	PALETTE6:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1:0]} == 6'b110111)	?	PALETTE7:
// Hires GR
// 2 color
			({COCO,BP,CRES,CHAR_LATCH[4]} == 5'b01000)							?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[4]} == 5'b01001)							?	PALETTE1:
// 4 Color
			({COCO,BP,CRES,ATRIB_LATCH[1:0]} == 6'b010100)						?	PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[1:0]} == 6'b010101)						?	PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH[1:0]} == 6'b010110)						?	PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH[1:0]} == 6'b010111)						?	PALETTE3:
// 16 color
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01100000)						?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01100001)						?	PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01100010)						?	PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01100011)						?	PALETTE3:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01100100)						?	PALETTE4:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01100101)						?	PALETTE5:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01100110)						?	PALETTE6:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01100111)						?	PALETTE7:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01101000)						?	PALETTE8:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01101001)						?	PALETTE9:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01101010)						?	PALETTEA:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01101011)						?	PALETTEB:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01101100)						?	PALETTEC:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01101101)						?	PALETTED:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01101110)						?	PALETTEE:
			({COCO,BP,CRES,CHAR_LATCH3[3:0]} == 8'b01101111)						?	PALETTEF:
																									PALETTE0;

assign PIXEL5 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,CHAR_LATCH[7],CHARACTER1[5]} == 6'b100001)			?	PALETTEC:
			({COCO,V,CHAR_LATCH[7],CHARACTER1[5]} == 6'b100000)			?	PALETTED:
// HR Text 80 (2 bytes is 1-8 pixel character)
// HR Text 40 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[5:3]}==7'b0011000)	?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[5:3]}==7'b0011001)	?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[5:3]}==7'b0011010)	?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[5:3]}==7'b0011011)	?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[5:3]}==7'b0011100)	?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[5:3]}==7'b0011101)	?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[5:3]}==7'b0011110)	?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[5:3]}==7'b0011111)	?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[2:0]}==7'b0010000)	?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[2:0]}==7'b0010001)	?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[2:0]}==7'b0010010)	?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[2:0]}==7'b0010011)	?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[2:0]}==7'b0010100)	?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[2:0]}==7'b0010101)	?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[2:0]}==7'b0010110)	?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER1[5],ATRIB_LATCH[2:0]}==7'b0010111)	?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER1[5]}==4'b0001)							?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[5]}==4'b0000)							?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[5]} == 5'b11111) ? PALETTEB:
// 4 COLOR
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3:2]} == 6'b110000)	?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3:2]} == 6'b110001)	?	PALETTE1:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3:2]} == 6'b110010)	?	PALETTE2:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3:2]} == 6'b110011)	?	PALETTE3:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3:2]} == 6'b110100)	?	PALETTE4:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3:2]} == 6'b110101)	?	PALETTE5:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3:2]} == 6'b110110)	?	PALETTE6:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3:2]} == 6'b110111)	?	PALETTE7:
// Hires GR
// 2 color
			({COCO,BP,CRES,CHAR_LATCH[5]} == 5'b01000)							?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[5]} == 5'b01001)							?	PALETTE1:
// 4 Color
			({COCO,BP,CRES,ATRIB_LATCH[3:2]} == 6'b010100)						?	PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[3:2]} == 6'b010101)						?	PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH[3:2]} == 6'b010110)						?	PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH[3:2]} == 6'b010111)						?	PALETTE3:
// 16 color
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01100000)						?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01100001)						?	PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01100010)						?	PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01100011)						?	PALETTE3:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01100100)						?	PALETTE4:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01100101)						?	PALETTE5:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01100110)						?	PALETTE6:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01100111)						?	PALETTE7:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01101000)						?	PALETTE8:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01101001)						?	PALETTE9:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01101010)						?	PALETTEA:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01101011)						?	PALETTEB:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01101100)						?	PALETTEC:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01101101)						?	PALETTED:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01101110)						?	PALETTEE:
			({COCO,BP,CRES,CHAR_LATCH3[7:4]} == 8'b01101111)						?	PALETTEF:
																									PALETTE0;

assign PIXEL6 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,CHAR_LATCH[7],CHARACTER1[6]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,CHAR_LATCH[7],CHARACTER1[6]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR Text 80 (2 bytes is 1-8 pixel character)
// HR Text 40 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER1[6],ATRIB_LATCH[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER1[6]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[6]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[6]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[6]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[6]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[6]} == 5'b11111) ? PALETTEB:
// 4 COLOR
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5:4]} == 6'b110000)	?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5:4]} == 6'b110001)	?	PALETTE1:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5:4]} == 6'b110010)	?	PALETTE2:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5:4]} == 6'b110011)	?	PALETTE3:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5:4]} == 6'b110100)	?	PALETTE4:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5:4]} == 6'b110101)	?	PALETTE5:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5:4]} == 6'b110110)	?	PALETTE6:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5:4]} == 6'b110111)	?	PALETTE7:
// Hires GR
// 2 color
			({COCO,BP,CRES,CHAR_LATCH[6]} == 5'b01000)							?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[6]} == 5'b01001)							?	PALETTE1:
// 4 Color
			({COCO,BP,CRES,ATRIB_LATCH[5:4]} == 6'b010100)						?	PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[5:4]} == 6'b010101)						?	PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH[5:4]} == 6'b010110)						?	PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH[5:4]} == 6'b010111)						?	PALETTE3:
// 16 color
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01100000)						?	PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01100001)						?	PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01100010)						?	PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01100011)						?	PALETTE3:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01100100)						?	PALETTE4:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01100101)						?	PALETTE5:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01100110)						?	PALETTE6:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01100111)						?	PALETTE7:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01101000)						?	PALETTE8:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01101001)						?	PALETTE9:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01101010)						?	PALETTEA:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01101011)						?	PALETTEB:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01101100)						?	PALETTEC:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01101101)						?	PALETTED:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01101110)						?	PALETTEE:
			({COCO,BP,CRES,ATRIB_LATCH3[3:0]} == 8'b01101111)						?	PALETTEF:
																									PALETTE0;

assign PIXEL7 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,CHAR_LATCH[7],CHARACTER1[7]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,CHAR_LATCH[7],CHARACTER1[7]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR Text 80 (2 bytes is 1-8 pixel character)
// HR Text 40 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER1[7],ATRIB_LATCH[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER1[7]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER1[7]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,CHAR_LATCH[7]} == 5'b11111) ? PALETTEB:
// 4 COLOR
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7:6]} == 6'b110000)	?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7:6]} == 6'b110001)	?	PALETTE1:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7:6]} == 6'b110010)	?	PALETTE2:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7:6]} == 6'b110011)	?	PALETTE3:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7:6]} == 6'b110100)	?	PALETTE4:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7:6]} == 6'b110101)	?	PALETTE5:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7:6]} == 6'b110110)	?	PALETTE6:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7:6]} == 6'b110111)	?	PALETTE7:
// Hires GR
// 2 color
			({COCO,BP,CRES,CHAR_LATCH[7]} == 5'b01000)							?	PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH[7]} == 5'b01001)							?	PALETTE1:
// 4 Color
			({COCO,BP,CRES,ATRIB_LATCH[7:6]} == 6'b010100)						?	PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[7:6]} == 6'b010101)						?	PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH[7:6]} == 6'b010110)						?	PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH[7:6]} == 6'b010111)						?	PALETTE3:
// 16 color
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01100000)						?	PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01100001)						?	PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01100010)						?	PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01100011)						?	PALETTE3:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01100100)						?	PALETTE4:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01100101)						?	PALETTE5:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01100110)						?	PALETTE6:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01100111)						?	PALETTE7:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01101000)						?	PALETTE8:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01101001)						?	PALETTE9:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01101010)						?	PALETTEA:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01101011)						?	PALETTEB:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01101100)						?	PALETTEC:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01101101)						?	PALETTED:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01101110)						?	PALETTEE:
			({COCO,BP,CRES,ATRIB_LATCH3[7:4]} == 8'b01101111)						?	PALETTEF:
																									PALETTE0;

assign PIXEL8 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[0]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[0]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR Text 80 (2 bytes is 1-8 pixel character)
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER3[0],ATRIB_LATCH3[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER4[0]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER4[0]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[0]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[0]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[0]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[0]} == 5'b11111) ? PALETTEB:
// Hires GR
// 2 color
			({COCO,BP,CRES,ATRIB_LATCH[0]} == 5'b01000) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[0]} == 5'b01001) ? PALETTE1:
// 4 Color
			({COCO,BP,CRES,CHAR_LATCH3[1:0]} == 6'b010100) ? PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH3[1:0]} == 6'b010101) ? PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH3[1:0]} == 6'b010110) ? PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH3[1:0]} == 6'b010111) ? PALETTE3:
																									PALETTE0;

assign PIXEL9 =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[1]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[1]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR text 80
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER3[1],ATRIB_LATCH3[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER4[1]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER4[1]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[1]} == 5'b11111) ? PALETTEB:
// Hires GR
// 2 color
			({COCO,BP,CRES,ATRIB_LATCH[1]} == 5'b01000) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[1]} == 5'b01001) ? PALETTE1:
// 4 Color
			({COCO,BP,CRES,CHAR_LATCH3[3:2]} == 6'b010100) ? PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH3[3:2]} == 6'b010101) ? PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH3[3:2]} == 6'b010110) ? PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH3[3:2]} == 6'b010111) ? PALETTE3:
																									PALETTE0;

assign PIXELA =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[2]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[2]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR text 80
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER3[2],ATRIB_LATCH3[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER4[2]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER4[2]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[2]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[2]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[2]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[2]} == 5'b11111) ? PALETTEB:
// Hires GR
// 2 color
			({COCO,BP,CRES,ATRIB_LATCH[2]} == 5'b01000) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[2]} == 5'b01001) ? PALETTE1:
// 4 Color
			({COCO,BP,CRES,CHAR_LATCH3[5:4]} == 6'b010100) ? PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH3[5:4]} == 6'b010101) ? PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH3[5:4]} == 6'b010110) ? PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH3[5:4]} == 6'b010111) ? PALETTE3:
																									PALETTE0;

assign PIXELB =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[3]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[3]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR text 80
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER3[3],ATRIB_LATCH3[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER4[3]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER4[3]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[3]} == 5'b11111) ? PALETTEB:
// Hires GR
// 2 color
			({COCO,BP,CRES,ATRIB_LATCH[3]} == 5'b01000) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[3]} == 5'b01001) ? PALETTE1:
// 4 Color
			({COCO,BP,CRES,CHAR_LATCH3[7:6]} == 6'b010100) ? PALETTE0:
			({COCO,BP,CRES,CHAR_LATCH3[7:6]} == 6'b010101) ? PALETTE1:
			({COCO,BP,CRES,CHAR_LATCH3[7:6]} == 6'b010110) ? PALETTE2:
			({COCO,BP,CRES,CHAR_LATCH3[7:6]} == 6'b010111) ? PALETTE3:
																									PALETTE0;

assign PIXELC =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[4]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[4]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR text 80
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER3[4],ATRIB_LATCH3[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER4[4]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER4[4]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[4]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[4]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[4]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[4]} == 5'b11111) ? PALETTEB:
// Hires GR
// 2 color
			({COCO,BP,CRES,ATRIB_LATCH[4]} == 5'b01000) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[4]} == 5'b01001) ? PALETTE1:
// 4 Color
			({COCO,BP,CRES,ATRIB_LATCH3[1:0]} == 6'b010100) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH3[1:0]} == 6'b010101) ? PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH3[1:0]} == 6'b010110) ? PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH3[1:0]} == 6'b010111) ? PALETTE3:
																									PALETTE0;

assign PIXELD =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[5]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[5]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR text 80
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER3[5],ATRIB_LATCH3[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER4[5]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER4[5]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[5]} == 5'b11111) ? PALETTEB:
// Hires GR
// 2 color
			({COCO,BP,CRES,ATRIB_LATCH[5]} == 5'b01000) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[5]} == 5'b01001) ? PALETTE1:
// 4 Color
			({COCO,BP,CRES,ATRIB_LATCH3[3:2]} == 6'b010100) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH3[3:2]} == 6'b010101) ? PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH3[3:2]} == 6'b010110) ? PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH3[3:2]} == 6'b010111) ? PALETTE3:
																									PALETTE0;

assign PIXELE =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[6]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[6]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR text 80
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER3[6],ATRIB_LATCH3[2:0]}==7'b0010111)?	PALETTE7:
// XTEXT 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER4[6]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER4[6]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[6]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[6]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[6]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[6]} == 5'b11111) ? PALETTEB:
// Hires GR
// 2 color
			({COCO,BP,CRES,ATRIB_LATCH[6]} == 5'b01000) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[6]} == 5'b01001) ? PALETTE1:
// 4 Color
			({COCO,BP,CRES,ATRIB_LATCH3[5:4]} == 6'b010100) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH3[5:4]} == 6'b010101) ? PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH3[5:4]} == 6'b010110) ? PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH3[5:4]} == 6'b010111) ? PALETTE3:
																									PALETTE0;

assign PIXELF =
//CoCo1 Text (2 bytes is 2-8 pixel characters) First byte
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[7]} == 6'b100001)	?	PALETTEC:		// Text On Inverted
			({COCO,V,ATRIB_LATCH[7],CHARACTER4[7]} == 6'b100000)	?	PALETTED:		// Text Off Inverted
// HR text 80
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[5:3]}==7'b0011000)?	PALETTE8:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[5:3]}==7'b0011001)?	PALETTE9:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[5:3]}==7'b0011010)?	PALETTEA:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[5:3]}==7'b0011011)?	PALETTEB:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[5:3]}==7'b0011100)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[5:3]}==7'b0011101)?	PALETTED:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[5:3]}==7'b0011110)?	PALETTEE:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[5:3]}==7'b0011111)?	PALETTEF:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[2:0]}==7'b0010000)?	PALETTE0:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[2:0]}==7'b0010001)?	PALETTE1:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[2:0]}==7'b0010010)?	PALETTE2:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[2:0]}==7'b0010011)?	PALETTE3:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[2:0]}==7'b0010100)?	PALETTE4:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[2:0]}==7'b0010101)?	PALETTE5:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[2:0]}==7'b0010110)?	PALETTE6:
			({COCO,BP,CRES[0],CHARACTER3[7],ATRIB_LATCH3[2:0]}==7'b0010111)?	PALETTE7:
// Lores 40 and 80 (2 bytes is 2-8 pixel characters)
			({COCO,BP,CRES[0],CHARACTER4[7]}==4'b0001)?	PALETTEC:
			({COCO,BP,CRES[0],CHARACTER4[7]}==4'b0000)?	PALETTED:
// Lowres graphics
// 2 color
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7]} == 5'b11100) ? PALETTE8:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7]} == 5'b11101) ? PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7]} == 5'b11110) ? PALETTEA:
			({COCO,COCO_GR,VID_CONT[0],CSS,ATRIB_LATCH[7]} == 5'b11111) ? PALETTEB:
// Hires GR
// 2 color
			({COCO,BP,CRES,ATRIB_LATCH[7]} == 5'b01000) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH[7]} == 5'b01001) ? PALETTE1:
// 4 Color
			({COCO,BP,CRES,ATRIB_LATCH3[7:6]} == 6'b010100) ? PALETTE0:
			({COCO,BP,CRES,ATRIB_LATCH3[7:6]} == 6'b010101) ? PALETTE1:
			({COCO,BP,CRES,ATRIB_LATCH3[7:6]} == 6'b010110) ? PALETTE2:
			({COCO,BP,CRES,ATRIB_LATCH3[7:6]} == 6'b010111) ? PALETTE3:
																									PALETTE0;

/*****************************************************************************
* Generate RGB
******************************************************************************/
// coco1 char		4:1		for 32 total pixels / 16 total pixels per byte / 8 pixels per byte
// coco3	40/no		4:1		for 32 total pixels / 16 pixels per byte
//	coco3 80/no		3:0		for 16 total pixels / 8 pixels per byte

// coco3 40/w		3:1		for 16 total pixels / 4 pixels per byte
// coco3 80/w		2:0		for 8 total pixels / 8 pixels per byte

assign PIXEL_ORDER =
// CoCo1 Text
// We display the after 16 bits so PIXEL_COUNT[4] needs to be inverted
							({COCO,COCO_GR,PIXEL_COUNT[4], CHAR_LATCH[7]} == 4'b1000)		?	4'b0000: // first 8 into 16 pixels
							({COCO,COCO_GR,PIXEL_COUNT[4],ATRIB_LATCH[7]} == 4'b1010)		?	4'b0001: // second 8 into 16 pixels
//	HR Text
// 32 / 40
							({COCO,BP,HRES[2],CRES[0]} == 4'b0001)									?	4'b0000:	// 32 / 40
// 64 / 80
							({COCO,BP,HRES[2],CRES[0]} == 4'b0011)									?	4'b0010:	//64 / 80
// XTEXT
// 32 / 40
							({COCO,BP,HRES[2],CRES[0],PIXEL_COUNT[4]} == 5'b00000)			?	4'b0000:	// 32 / 40
							({COCO,BP,HRES[2],CRES[0],PIXEL_COUNT[4]} == 5'b00001)			?	4'b0001:	// 32 / 40
// 64 / 80
							({COCO,BP,HRES[2],CRES[0]} == 4'b0010)									?	4'b0011:	//64 / 80
// SG4
							({COCO,COCO_GR,PIXEL_COUNT[4], CHAR_LATCH[7]} == 4'b1001)		?	4'b1001:
							({COCO,COCO_GR,PIXEL_COUNT[4],ATRIB_LATCH[7]} == 4'b1011)		?	4'b1000:
// Lowres graphics
// 256 2 identicle pixels in a row
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[4]} == 6'b111110)			?	4'b0000: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[4]} == 6'b111111)			?	4'b0001: // second 8 into 16 pixels
// 128x4 4 identicle pixels in a row
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[4]} == 6'b110100)			?	4'b0100: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[4]} == 6'b110101)			?	4'b0101: // second 8 into 16 pixels

							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[4]} == 6'b111000)			?	4'b0100: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[4]} == 6'b111001)			?	4'b0101: // second 8 into 16 pixels

							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[4]} == 6'b111100)			?	4'b0100: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[4]} == 6'b111101)			?	4'b0101: // second 8 into 16 pixels
// 128x2 4 identicle pixels in a row
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1100101)		?	4'b0100: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1100100)		?	4'b0101: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1100111)		?	4'b0110: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1100110)		?	4'b0111: // second 8 into 16 pixels

							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1101101)		?	4'b0100: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1101100)		?	4'b0101: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1101111)		?	4'b0110: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1101110)		?	4'b0111: // second 8 into 16 pixels

							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1110101)		?	4'b0100: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1110100)		?	4'b0101: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1110111)		?	4'b0110: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1110110)		?	4'b0111: // second 8 into 16 pixels
// 64 8 identicle pixels in a row
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1100001)		?	4'b1000: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1100000)		?	4'b1001: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1100011)		?	4'b1010: // second 8 into 16 pixels
							({COCO,COCO_GR,VID_CONT[2:0],PIXEL_COUNT[5:4]} == 7'b1100010)		?	4'b1011: // second 8 into 16 pixels
// HR GR
// 512X4
							({COCO,BP,HRES[2:1],CRES} == 6'b011101)									?	4'b1100:
// 512X2
							({COCO,BP,HRES[2:1],CRES} == 6'b011000)									?	4'b1010:
// 256x16
							({COCO,BP,HRES[2:1],CRES} == 6'b011110)									?	4'b1110:
// 256X4
							({COCO,BP,HRES[2:1],CRES} == 6'b011001)								 	?	4'b1011:
// 256X2
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[4]} == 7'b0101000)				?	4'b0000:
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[4]} == 7'b0101001)				?	4'b0001:
// 128x16
							({COCO,BP,HRES[2:1],CRES} == 6'b011010)									?	4'b1101:
// 128X4
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[4]} == 7'b0101010)				?	4'b0100:
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[4]} == 7'b0101011)				?	4'b0101:
// 128X2
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[5:4]} == 8'b01000000)			?	4'b0100:
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[5:4]} == 8'b01000001)			?	4'b0101:
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[5:4]} == 8'b01000010)			?	4'b0110:
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[5:4]} == 8'b01000011)			?	4'b0111:
// 64X16
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[4]} == 7'b0100100)				?	4'b1000:
							({COCO,BP,HRES[2:1],CRES,PIXEL_COUNT[4]} == 7'b0100101)				?	4'b1001:

																														4'b0000;

always @ (negedge PIX_CLK)
begin
	RED1 <= RED1X;
	GREEN1 <= GREEN1X;
	BLUE1 <= BLUE1X;
	RED0 <= RED0X;
	GREEN0 <= GREEN0X;
	BLUE0 <= BLUE0X;
	if(PIXEL_COUNT[3:0] == 4'b1111)
	begin
		case (PIXEL_ORDER)
		default:	// 0x0000
		begin
// Displayed pixels mare 2x real pixels first half
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL7[5],PIXEL7[5],PIXEL6[5],PIXEL6[5],PIXEL5[5],PIXEL5[5],PIXEL4[5],PIXEL4[5],PIXEL3[5],PIXEL3[5],PIXEL2[5],PIXEL2[5],PIXEL1[5],PIXEL1[5],PIXEL0[5],PIXEL0[5]};
			GREEN1S <=	{PIXEL7[4],PIXEL7[4],PIXEL6[4],PIXEL6[4],PIXEL5[4],PIXEL5[4],PIXEL4[4],PIXEL4[4],PIXEL3[4],PIXEL3[4],PIXEL2[4],PIXEL2[4],PIXEL1[4],PIXEL1[4],PIXEL0[4],PIXEL0[4]};
			BLUE1S <=	{PIXEL7[3],PIXEL7[3],PIXEL6[3],PIXEL6[3],PIXEL5[3],PIXEL5[3],PIXEL4[3],PIXEL4[3],PIXEL3[3],PIXEL3[3],PIXEL2[3],PIXEL2[3],PIXEL1[3],PIXEL1[3],PIXEL0[3],PIXEL0[3]};
			RED0S <=		{PIXEL7[2],PIXEL7[2],PIXEL6[2],PIXEL6[2],PIXEL5[2],PIXEL5[2],PIXEL4[2],PIXEL4[2],PIXEL3[2],PIXEL3[2],PIXEL2[2],PIXEL2[2],PIXEL1[2],PIXEL1[2],PIXEL0[2],PIXEL0[2]};
			GREEN0S <=	{PIXEL7[1],PIXEL7[1],PIXEL6[1],PIXEL6[1],PIXEL5[1],PIXEL5[1],PIXEL4[1],PIXEL4[1],PIXEL3[1],PIXEL3[1],PIXEL2[1],PIXEL2[1],PIXEL1[1],PIXEL1[1],PIXEL0[1],PIXEL0[1]};
			BLUE0S <=	{PIXEL7[0],PIXEL7[0],PIXEL6[0],PIXEL6[0],PIXEL5[0],PIXEL5[0],PIXEL4[0],PIXEL4[0],PIXEL3[0],PIXEL3[0],PIXEL2[0],PIXEL2[0],PIXEL1[0],PIXEL1[0],PIXEL0[0],PIXEL0[0]};
		end
		4'b0001:
		begin
// Displayed pixels mare 2x real pixels second half
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXELF[5],PIXELF[5],PIXELE[5],PIXELE[5],PIXELD[5],PIXELD[5],PIXELC[5],PIXELC[5],PIXELB[5],PIXELB[5],PIXELA[5],PIXELA[5],PIXEL9[5],PIXEL9[5],PIXEL8[5],PIXEL8[5]};
			GREEN1S <=	{PIXELF[4],PIXELF[4],PIXELE[4],PIXELE[4],PIXELD[4],PIXELD[4],PIXELC[4],PIXELC[4],PIXELB[4],PIXELB[4],PIXELA[4],PIXELA[4],PIXEL9[4],PIXEL9[4],PIXEL8[4],PIXEL8[4]};
			BLUE1S <=	{PIXELF[3],PIXELF[3],PIXELE[3],PIXELE[3],PIXELD[3],PIXELD[3],PIXELC[3],PIXELC[3],PIXELB[3],PIXELB[3],PIXELA[3],PIXELA[3],PIXEL9[3],PIXEL9[3],PIXEL8[3],PIXEL8[3]};
			RED0S <=		{PIXELF[2],PIXELF[2],PIXELE[2],PIXELE[2],PIXELD[2],PIXELD[2],PIXELC[2],PIXELC[2],PIXELB[2],PIXELB[2],PIXELA[2],PIXELA[2],PIXEL9[2],PIXEL9[2],PIXEL8[2],PIXEL8[2]};
			GREEN0S <=	{PIXELF[1],PIXELF[1],PIXELE[1],PIXELE[1],PIXELD[1],PIXELD[1],PIXELC[1],PIXELC[1],PIXELB[1],PIXELB[1],PIXELA[1],PIXELA[1],PIXEL9[1],PIXEL9[1],PIXEL8[1],PIXEL8[1]};
			BLUE0S <=	{PIXELF[0],PIXELF[0],PIXELE[0],PIXELE[0],PIXELD[0],PIXELD[0],PIXELC[0],PIXELC[0],PIXELB[0],PIXELB[0],PIXELA[0],PIXELA[0],PIXEL9[0],PIXEL9[0],PIXEL8[0],PIXEL8[0]};
		end
		4'b0010:
		begin
// Displayed pixels are 1x
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXELF[5],PIXELE[5],PIXELD[5],PIXELC[5],PIXELB[5],PIXELA[5],PIXEL9[5],PIXEL8[5],PIXEL7[5],PIXEL6[5],PIXEL5[5],PIXEL4[5],PIXEL3[5],PIXEL2[5],PIXEL1[5],PIXEL0[5]};
			GREEN1S <=	{PIXELF[4],PIXELE[4],PIXELD[4],PIXELC[4],PIXELB[4],PIXELA[4],PIXEL9[4],PIXEL8[4],PIXEL7[4],PIXEL6[4],PIXEL5[4],PIXEL4[4],PIXEL3[4],PIXEL2[4],PIXEL1[4],PIXEL0[4]};
			BLUE1S <=	{PIXELF[3],PIXELE[3],PIXELD[3],PIXELC[3],PIXELB[3],PIXELA[3],PIXEL9[3],PIXEL8[3],PIXEL7[3],PIXEL6[3],PIXEL5[3],PIXEL4[3],PIXEL3[3],PIXEL2[3],PIXEL1[3],PIXEL0[3]};
			RED0S <=		{PIXELF[2],PIXELE[2],PIXELD[2],PIXELC[2],PIXELB[2],PIXELA[2],PIXEL9[2],PIXEL8[2],PIXEL7[2],PIXEL6[2],PIXEL5[2],PIXEL4[2],PIXEL3[2],PIXEL2[2],PIXEL1[2],PIXEL0[2]};
			GREEN0S <=	{PIXELF[1],PIXELE[1],PIXELD[1],PIXELC[1],PIXELB[1],PIXELA[1],PIXEL9[1],PIXEL8[1],PIXEL7[1],PIXEL6[1],PIXEL5[1],PIXEL4[1],PIXEL3[1],PIXEL2[1],PIXEL1[1],PIXEL0[1]};
			BLUE0S <=	{PIXELF[0],PIXELE[0],PIXELD[0],PIXELC[0],PIXELB[0],PIXELA[0],PIXEL9[0],PIXEL8[0],PIXEL7[0],PIXEL6[0],PIXEL5[0],PIXEL4[0],PIXEL3[0],PIXEL2[0],PIXEL1[0],PIXEL0[0]};
		end
		4'b0011:
		begin
// Displayed pixels are 1x
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL7[5],PIXEL6[5],PIXEL5[5],PIXEL4[5],PIXEL3[5],PIXEL2[5],PIXEL1[5],PIXEL0[5],PIXELF[5],PIXELE[5],PIXELD[5],PIXELC[5],PIXELB[5],PIXELA[5],PIXEL9[5],PIXEL8[5]};
			GREEN1S <=	{PIXEL7[4],PIXEL6[4],PIXEL5[4],PIXEL4[4],PIXEL3[4],PIXEL2[4],PIXEL1[4],PIXEL0[4],PIXELF[4],PIXELE[4],PIXELD[4],PIXELC[4],PIXELB[4],PIXELA[4],PIXEL9[4],PIXEL8[4]};
			BLUE1S <=	{PIXEL7[3],PIXEL6[3],PIXEL5[3],PIXEL4[3],PIXEL3[3],PIXEL2[3],PIXEL1[3],PIXEL0[3],PIXELF[3],PIXELE[3],PIXELD[3],PIXELC[3],PIXELB[3],PIXELA[3],PIXEL9[3],PIXEL8[3]};
			RED0S <=		{PIXEL7[2],PIXEL6[2],PIXEL5[2],PIXEL4[2],PIXEL3[2],PIXEL2[2],PIXEL1[2],PIXEL0[2],PIXELF[2],PIXELE[2],PIXELD[2],PIXELC[2],PIXELB[2],PIXELA[2],PIXEL9[2],PIXEL8[2]};
			GREEN0S <=	{PIXEL7[1],PIXEL6[1],PIXEL5[1],PIXEL4[1],PIXEL3[1],PIXEL2[1],PIXEL1[1],PIXEL0[1],PIXELF[1],PIXELE[1],PIXELD[1],PIXELC[1],PIXELB[1],PIXELA[1],PIXEL9[1],PIXEL8[1]};
			BLUE0S <=	{PIXEL7[0],PIXEL6[0],PIXEL5[0],PIXEL4[0],PIXEL3[0],PIXEL2[0],PIXEL1[0],PIXEL0[0],PIXELF[0],PIXELE[0],PIXELD[0],PIXELC[0],PIXELB[0],PIXELA[0],PIXEL9[0],PIXEL8[0]};
		end
		4'b0100:
		begin
// Displayed pixels are 4x real pixels
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL2[5],PIXEL2[5],PIXEL2[5],PIXEL2[5],PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL0[5],PIXEL0[5],PIXEL0[5],PIXEL0[5]};
			GREEN1S <=	{PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL2[4],PIXEL2[4],PIXEL2[4],PIXEL2[4],PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL0[4],PIXEL0[4],PIXEL0[4],PIXEL0[4]};
			BLUE1S <=	{PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL2[3],PIXEL2[3],PIXEL2[3],PIXEL2[3],PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL0[3],PIXEL0[3],PIXEL0[3],PIXEL0[3]};
			RED0S <=		{PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL2[2],PIXEL2[2],PIXEL2[2],PIXEL2[2],PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL0[2],PIXEL0[2],PIXEL0[2],PIXEL0[2]};
			GREEN0S <=	{PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL2[1],PIXEL2[1],PIXEL2[1],PIXEL2[1],PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL0[1],PIXEL0[1],PIXEL0[1],PIXEL0[1]};
			BLUE0S <=	{PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL2[0],PIXEL2[0],PIXEL2[0],PIXEL2[0],PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL0[0],PIXEL0[0],PIXEL0[0],PIXEL0[0]};
		end
		4'b0101:
		begin
// Displayed pixels are 4x reaL pixels
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL7[5],PIXEL7[5],PIXEL7[5],PIXEL7[5],PIXEL6[5],PIXEL6[5],PIXEL6[5],PIXEL6[5],PIXEL5[5],PIXEL5[5],PIXEL5[5],PIXEL5[5],PIXEL4[5],PIXEL4[5],PIXEL4[5],PIXEL4[5]};
			GREEN1S <=	{PIXEL7[4],PIXEL7[4],PIXEL7[4],PIXEL7[4],PIXEL6[4],PIXEL6[4],PIXEL6[4],PIXEL6[4],PIXEL5[4],PIXEL5[4],PIXEL5[4],PIXEL5[4],PIXEL4[4],PIXEL4[4],PIXEL4[4],PIXEL4[4]};
			BLUE1S <=	{PIXEL7[3],PIXEL7[3],PIXEL7[3],PIXEL7[3],PIXEL6[3],PIXEL6[3],PIXEL6[3],PIXEL6[3],PIXEL5[3],PIXEL5[3],PIXEL5[3],PIXEL5[3],PIXEL4[3],PIXEL4[3],PIXEL4[3],PIXEL4[3]};
			RED0S <=		{PIXEL7[2],PIXEL7[2],PIXEL7[2],PIXEL7[2],PIXEL6[2],PIXEL6[2],PIXEL6[2],PIXEL6[2],PIXEL5[2],PIXEL5[2],PIXEL5[2],PIXEL5[2],PIXEL4[2],PIXEL4[2],PIXEL4[2],PIXEL4[2]};
			GREEN0S <=	{PIXEL7[1],PIXEL7[1],PIXEL7[1],PIXEL7[1],PIXEL6[1],PIXEL6[1],PIXEL6[1],PIXEL6[1],PIXEL5[1],PIXEL5[1],PIXEL5[1],PIXEL5[1],PIXEL4[1],PIXEL4[1],PIXEL4[1],PIXEL4[1]};
			BLUE0S <=	{PIXEL7[0],PIXEL7[0],PIXEL7[0],PIXEL7[0],PIXEL6[0],PIXEL6[0],PIXEL6[0],PIXEL6[0],PIXEL5[0],PIXEL5[0],PIXEL5[0],PIXEL5[0],PIXEL4[0],PIXEL4[0],PIXEL4[0],PIXEL4[0]};
		end
		4'b0110:
		begin
// Displayed pixels are 4x real pixels
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXELB[5],PIXELB[5],PIXELB[5],PIXELB[5],PIXELA[5],PIXELA[5],PIXELA[5],PIXELA[5],PIXEL9[5],PIXEL9[5],PIXEL9[5],PIXEL9[5],PIXEL8[5],PIXEL8[5],PIXEL8[5],PIXEL8[5]};
			GREEN1S <=	{PIXELB[4],PIXELB[4],PIXELB[4],PIXELB[4],PIXELA[4],PIXELA[4],PIXELA[4],PIXELA[4],PIXEL9[4],PIXEL9[4],PIXEL9[4],PIXEL9[4],PIXEL8[4],PIXEL8[4],PIXEL8[4],PIXEL8[4]};
			BLUE1S <=	{PIXELB[3],PIXELB[3],PIXELB[3],PIXELB[3],PIXELA[3],PIXELA[3],PIXELA[3],PIXELA[3],PIXEL9[3],PIXEL9[3],PIXEL9[3],PIXEL9[3],PIXEL8[3],PIXEL8[3],PIXEL8[3],PIXEL8[3]};
			RED0S <=		{PIXELB[2],PIXELB[2],PIXELB[2],PIXELB[2],PIXELA[2],PIXELA[2],PIXELA[2],PIXELA[2],PIXEL9[2],PIXEL9[2],PIXEL9[2],PIXEL9[2],PIXEL8[2],PIXEL8[2],PIXEL8[2],PIXEL8[2]};
			GREEN0S <=	{PIXELB[1],PIXELB[1],PIXELB[1],PIXELB[1],PIXELA[1],PIXELA[1],PIXELA[1],PIXELA[1],PIXEL9[1],PIXEL9[1],PIXEL9[1],PIXEL9[1],PIXEL8[1],PIXEL8[1],PIXEL8[1],PIXEL8[1]};
			BLUE0S <=	{PIXELB[0],PIXELB[0],PIXELB[0],PIXELB[0],PIXELA[0],PIXELA[0],PIXELA[0],PIXELA[0],PIXEL9[0],PIXEL9[0],PIXEL9[0],PIXEL9[0],PIXEL8[0],PIXEL8[0],PIXEL8[0],PIXEL8[0]};
		end
		4'b0111:
		begin
// Displayed pixels are 4x real pixelS
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXELF[5],PIXELF[5],PIXELF[5],PIXELF[5],PIXELE[5],PIXELE[5],PIXELE[5],PIXELE[5],PIXELD[5],PIXELD[5],PIXELD[5],PIXELD[5],PIXELC[5],PIXELC[5],PIXELC[5],PIXELC[5]};
			GREEN1S <=	{PIXELF[4],PIXELF[4],PIXELF[4],PIXELF[4],PIXELE[4],PIXELE[4],PIXELE[4],PIXELE[4],PIXELD[4],PIXELD[4],PIXELD[4],PIXELD[4],PIXELC[4],PIXELC[4],PIXELC[4],PIXELC[4]};
			BLUE1S <=	{PIXELF[3],PIXELF[3],PIXELF[3],PIXELF[3],PIXELE[3],PIXELE[3],PIXELE[3],PIXELE[3],PIXELD[3],PIXELD[3],PIXELD[3],PIXELD[3],PIXELC[3],PIXELC[3],PIXELC[3],PIXELC[3]};
			RED0S <=		{PIXELF[2],PIXELF[2],PIXELF[2],PIXELF[2],PIXELE[2],PIXELE[2],PIXELE[2],PIXELE[2],PIXELD[2],PIXELD[2],PIXELD[2],PIXELD[2],PIXELC[2],PIXELC[2],PIXELC[2],PIXELC[2]};
			GREEN0S <=	{PIXELF[1],PIXELF[1],PIXELF[1],PIXELF[1],PIXELE[1],PIXELE[1],PIXELE[1],PIXELE[1],PIXELD[1],PIXELD[1],PIXELD[1],PIXELD[1],PIXELC[1],PIXELC[1],PIXELC[1],PIXELC[1]};
			BLUE0S <=	{PIXELF[0],PIXELF[0],PIXELF[0],PIXELF[0],PIXELE[0],PIXELE[0],PIXELE[0],PIXELE[0],PIXELD[0],PIXELD[0],PIXELD[0],PIXELD[0],PIXELC[0],PIXELC[0],PIXELC[0],PIXELC[0]};
		end
		4'b1000:
		begin
// Displayed pixels mare 8x real pixels
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL2[5],PIXEL2[5],PIXEL2[5],PIXEL2[5],PIXEL2[5],PIXEL2[5],PIXEL2[5],PIXEL2[5]};
			GREEN1S <=	{PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL2[4],PIXEL2[4],PIXEL2[4],PIXEL2[4],PIXEL2[4],PIXEL2[4],PIXEL2[4],PIXEL2[4]};
			BLUE1S <=	{PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL2[3],PIXEL2[3],PIXEL2[3],PIXEL2[3],PIXEL2[3],PIXEL2[3],PIXEL2[3],PIXEL2[3]};
			RED0S <=		{PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL2[2],PIXEL2[2],PIXEL2[2],PIXEL2[2],PIXEL2[2],PIXEL2[2],PIXEL2[2],PIXEL2[2]};
			GREEN0S <=	{PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL2[1],PIXEL2[1],PIXEL2[1],PIXEL2[1],PIXEL2[1],PIXEL2[1],PIXEL2[1],PIXEL2[1]};
			BLUE0S <=	{PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL2[0],PIXEL2[0],PIXEL2[0],PIXEL2[0],PIXEL2[0],PIXEL2[0],PIXEL2[0],PIXEL2[0]};
		end
		4'b1001:
		begin
// Displayed pixels are 8x real pixels
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL0[5],PIXEL0[5],PIXEL0[5],PIXEL0[5],PIXEL0[5],PIXEL0[5],PIXEL0[5],PIXEL0[5]};
			GREEN1S <=	{PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL0[4],PIXEL0[4],PIXEL0[4],PIXEL0[4],PIXEL0[4],PIXEL0[4],PIXEL0[4],PIXEL0[4]};
			BLUE1S <=	{PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL0[3],PIXEL0[3],PIXEL0[3],PIXEL0[3],PIXEL0[3],PIXEL0[3],PIXEL0[3],PIXEL0[3]};
			RED0S <=		{PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL0[2],PIXEL0[2],PIXEL0[2],PIXEL0[2],PIXEL0[2],PIXEL0[2],PIXEL0[2],PIXEL0[2]};
			GREEN0S <=	{PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL0[1],PIXEL0[1],PIXEL0[1],PIXEL0[1],PIXEL0[1],PIXEL0[1],PIXEL0[1],PIXEL0[1]};
			BLUE0S <=	{PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL0[0],PIXEL0[0],PIXEL0[0],PIXEL0[0],PIXEL0[0],PIXEL0[0],PIXEL0[0],PIXEL0[0]};
		end
		4'b1010:
		begin
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL7[5],PIXEL6[5],PIXEL5[5],PIXEL4[5],PIXEL3[5],PIXEL2[5],PIXEL1[5],PIXEL0[5],PIXELF[5],PIXELE[5],PIXELD[5],PIXELC[5],PIXELB[5],PIXELA[5],PIXEL9[5],PIXEL8[5]};
			GREEN1S <=	{PIXEL7[4],PIXEL6[4],PIXEL5[4],PIXEL4[4],PIXEL3[4],PIXEL2[4],PIXEL1[4],PIXEL0[4],PIXELF[4],PIXELE[4],PIXELD[4],PIXELC[4],PIXELB[4],PIXELA[4],PIXEL9[4],PIXEL8[4]};
			BLUE1S <=	{PIXEL7[3],PIXEL6[3],PIXEL5[3],PIXEL4[3],PIXEL3[3],PIXEL2[3],PIXEL1[3],PIXEL0[3],PIXELF[3],PIXELE[3],PIXELD[3],PIXELC[3],PIXELB[3],PIXELA[3],PIXEL9[3],PIXEL8[3]};
			RED0S <=		{PIXEL7[2],PIXEL6[2],PIXEL5[2],PIXEL4[2],PIXEL3[2],PIXEL2[2],PIXEL1[2],PIXEL0[2],PIXELF[2],PIXELE[2],PIXELD[2],PIXELC[2],PIXELB[2],PIXELA[2],PIXEL9[2],PIXEL8[2]};
			GREEN0S <=	{PIXEL7[1],PIXEL6[1],PIXEL5[1],PIXEL4[1],PIXEL3[1],PIXEL2[1],PIXEL1[1],PIXEL0[1],PIXELF[1],PIXELE[1],PIXELD[1],PIXELC[1],PIXELB[1],PIXELA[1],PIXEL9[1],PIXEL8[1]};
			BLUE0S <=	{PIXEL7[0],PIXEL6[0],PIXEL5[0],PIXEL4[0],PIXEL3[0],PIXEL2[0],PIXEL1[0],PIXEL0[0],PIXELF[0],PIXELE[0],PIXELD[0],PIXELC[0],PIXELB[0],PIXELA[0],PIXEL9[0],PIXEL8[0]};
		end
		4'b1011:
		begin
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL3[5],PIXEL3[5],PIXEL2[5],PIXEL2[5],PIXEL1[5],PIXEL1[5],PIXEL0[5],PIXEL0[5],PIXEL7[5],PIXEL7[5],PIXEL6[5],PIXEL6[5],PIXEL5[5],PIXEL5[5],PIXEL4[5],PIXEL4[5]};
			GREEN1S <=	{PIXEL3[4],PIXEL3[4],PIXEL2[4],PIXEL2[4],PIXEL1[4],PIXEL1[4],PIXEL0[4],PIXEL0[4],PIXEL7[4],PIXEL7[4],PIXEL6[4],PIXEL6[4],PIXEL5[4],PIXEL5[4],PIXEL4[4],PIXEL4[4]};
			BLUE1S <=	{PIXEL3[3],PIXEL3[3],PIXEL2[3],PIXEL2[3],PIXEL1[3],PIXEL1[3],PIXEL0[3],PIXEL0[3],PIXEL7[3],PIXEL7[3],PIXEL6[3],PIXEL6[3],PIXEL5[3],PIXEL5[3],PIXEL4[3],PIXEL4[3]};
			RED0S <=		{PIXEL3[2],PIXEL3[2],PIXEL2[2],PIXEL2[2],PIXEL1[2],PIXEL1[2],PIXEL0[2],PIXEL0[2],PIXEL7[2],PIXEL7[2],PIXEL6[2],PIXEL6[2],PIXEL5[2],PIXEL5[2],PIXEL4[2],PIXEL4[2]};
			GREEN0S <=	{PIXEL3[1],PIXEL3[1],PIXEL2[1],PIXEL2[1],PIXEL1[1],PIXEL1[1],PIXEL0[1],PIXEL0[1],PIXEL7[1],PIXEL7[1],PIXEL6[1],PIXEL6[1],PIXEL5[1],PIXEL5[1],PIXEL4[1],PIXEL4[1]};
			BLUE0S <=	{PIXEL3[0],PIXEL3[0],PIXEL2[0],PIXEL2[0],PIXEL1[0],PIXEL1[0],PIXEL0[0],PIXEL0[0],PIXEL7[0],PIXEL7[0],PIXEL6[0],PIXEL6[0],PIXEL5[0],PIXEL5[0],PIXEL4[0],PIXEL4[0]};
		end
		4'b1100:
		begin
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXELB[5],PIXELA[5],PIXEL9[5],PIXEL8[5],PIXELF[5],PIXELE[5],PIXELD[5],PIXELC[5],PIXEL3[5],PIXEL2[5],PIXEL1[5],PIXEL0[5],PIXEL7[5],PIXEL6[5],PIXEL5[5],PIXEL4[5]};
			GREEN1S <=	{PIXELB[4],PIXELA[4],PIXEL9[4],PIXEL8[4],PIXELF[4],PIXELE[4],PIXELD[4],PIXELC[4],PIXEL3[4],PIXEL2[4],PIXEL1[4],PIXEL0[4],PIXEL7[4],PIXEL6[4],PIXEL5[4],PIXEL4[4]};
			BLUE1S <=	{PIXELB[3],PIXELA[3],PIXEL9[3],PIXEL8[3],PIXELF[3],PIXELE[3],PIXELD[3],PIXELC[3],PIXEL3[3],PIXEL2[3],PIXEL1[3],PIXEL0[3],PIXEL7[3],PIXEL6[3],PIXEL5[3],PIXEL4[3]};
			RED0S <=		{PIXELB[2],PIXELA[2],PIXEL9[2],PIXEL8[2],PIXELF[2],PIXELE[2],PIXELD[2],PIXELC[2],PIXEL3[2],PIXEL2[2],PIXEL1[2],PIXEL0[2],PIXEL7[2],PIXEL6[2],PIXEL5[2],PIXEL4[2]};
			GREEN0S <=	{PIXELB[1],PIXELA[1],PIXEL9[1],PIXEL8[1],PIXELF[1],PIXELE[1],PIXELD[1],PIXELC[1],PIXEL3[1],PIXEL2[1],PIXEL1[1],PIXEL0[1],PIXEL7[1],PIXEL6[1],PIXEL5[1],PIXEL4[1]};
			BLUE0S <=	{PIXELB[0],PIXELA[0],PIXEL9[0],PIXEL8[0],PIXELF[0],PIXELE[0],PIXELD[0],PIXELC[0],PIXEL3[0],PIXEL2[0],PIXEL1[0],PIXEL0[0],PIXEL7[0],PIXEL6[0],PIXEL5[0],PIXEL4[0]};
		end
		4'b1101:
		begin
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL1[5],PIXEL0[5],PIXEL0[5],PIXEL0[5],PIXEL0[5],PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL3[5],PIXEL2[5],PIXEL2[5],PIXEL2[5],PIXEL2[5]};
			GREEN1S <=	{PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL1[4],PIXEL0[4],PIXEL0[4],PIXEL0[4],PIXEL0[4],PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL3[4],PIXEL2[4],PIXEL2[4],PIXEL2[4],PIXEL2[4]};
			BLUE1S <=	{PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL1[3],PIXEL0[3],PIXEL0[3],PIXEL0[3],PIXEL0[3],PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL3[3],PIXEL2[3],PIXEL2[3],PIXEL2[3],PIXEL2[3]};
			RED0S <=		{PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL1[2],PIXEL0[2],PIXEL0[2],PIXEL0[2],PIXEL0[2],PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL3[2],PIXEL2[2],PIXEL2[2],PIXEL2[2],PIXEL2[2]};
			GREEN0S <=	{PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL1[1],PIXEL0[1],PIXEL0[1],PIXEL0[1],PIXEL0[1],PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL3[1],PIXEL2[1],PIXEL2[1],PIXEL2[1],PIXEL2[1]};
			BLUE0S <=	{PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL1[0],PIXEL0[0],PIXEL0[0],PIXEL0[0],PIXEL0[0],PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL3[0],PIXEL2[0],PIXEL2[0],PIXEL2[0],PIXEL2[0]};
		end
		4'b1110:
		begin
//                           15        14        13        12        11        10         9         8         7         6         5         4         3         2         1         0
			RED1S <=		{PIXEL5[5],PIXEL5[5],PIXEL4[5],PIXEL4[5],PIXEL7[5],PIXEL7[5],PIXEL6[5],PIXEL6[5],PIXEL1[5],PIXEL1[5],PIXEL0[5],PIXEL0[5],PIXEL3[5],PIXEL3[5],PIXEL2[5],PIXEL2[5]};
			GREEN1S <=	{PIXEL5[4],PIXEL5[4],PIXEL4[4],PIXEL4[4],PIXEL7[4],PIXEL7[4],PIXEL6[4],PIXEL6[4],PIXEL1[4],PIXEL1[4],PIXEL0[4],PIXEL0[4],PIXEL3[4],PIXEL3[4],PIXEL2[4],PIXEL2[4]};
			BLUE1S <=	{PIXEL5[3],PIXEL5[3],PIXEL4[3],PIXEL4[3],PIXEL7[3],PIXEL7[3],PIXEL6[3],PIXEL6[3],PIXEL1[3],PIXEL1[3],PIXEL0[3],PIXEL0[3],PIXEL3[3],PIXEL3[3],PIXEL2[3],PIXEL2[3]};
			RED0S <=		{PIXEL5[2],PIXEL5[2],PIXEL4[2],PIXEL4[2],PIXEL7[2],PIXEL7[2],PIXEL6[2],PIXEL6[2],PIXEL1[2],PIXEL1[2],PIXEL0[2],PIXEL0[2],PIXEL3[2],PIXEL3[2],PIXEL2[2],PIXEL2[2]};
			GREEN0S <=	{PIXEL5[1],PIXEL5[1],PIXEL4[1],PIXEL4[1],PIXEL7[1],PIXEL7[1],PIXEL6[1],PIXEL6[1],PIXEL1[1],PIXEL1[1],PIXEL0[1],PIXEL0[1],PIXEL3[1],PIXEL3[1],PIXEL2[1],PIXEL2[1]};
			BLUE0S <=	{PIXEL5[0],PIXEL5[0],PIXEL4[0],PIXEL4[0],PIXEL7[0],PIXEL7[0],PIXEL6[0],PIXEL6[0],PIXEL1[0],PIXEL1[0],PIXEL0[0],PIXEL0[0],PIXEL3[0],PIXEL3[0],PIXEL2[0],PIXEL2[0]};
		end
		endcase
	end
end

assign BORDER =
			({COCO,COCO_GR} == 2'b10)								?	6'b000000:
			({COCO,COCO_GR,VID_CONT[0],CSS} == 4'b1110)		?	PALETTE9:
			({COCO,COCO_GR,VID_CONT[0],CSS} == 4'b1111)		?	PALETTEB:
			({COCO,COCO_GR,VID_CONT[0],CSS} == 4'b1100)		?	PALETTE0:
			({COCO,COCO_GR,VID_CONT[0],CSS} == 4'b1101)		?	PALETTE4:
//COCO3
																				BDR_PAL;

assign RED1X =		({VBLANKING,HBLANKING} == 2'b00)				?	RED1S[~PIXEL_COUNT[3:0]]:
		({(VBORDER&HBORDER),(VBLANKING|HBLANKING)} == 2'b11)	?	BORDER[5]:
																					1'b0;

assign GREEN1X =	({VBLANKING,HBLANKING} == 2'b00)				?	GREEN1S[~PIXEL_COUNT[3:0]]:
		({(VBORDER&HBORDER),(VBLANKING|HBLANKING)} == 2'b11)	?	BORDER[4]:
																					1'b0;

assign BLUE1X =	({VBLANKING,HBLANKING} == 2'b00)				?	BLUE1S[~PIXEL_COUNT[3:0]]:
		({(VBORDER&HBORDER),(VBLANKING|HBLANKING)} == 2'b11)	?	BORDER[3]:
																					1'b0;

assign RED0X =		({VBLANKING,HBLANKING} == 2'b00)				?	RED0S[~PIXEL_COUNT[3:0]]:
		({(VBORDER&HBORDER),(VBLANKING|HBLANKING)} == 2'b11)	?	BORDER[2]:
																					1'b0;

assign GREEN0X =	({VBLANKING,HBLANKING} == 2'b00)				?	GREEN0S[~PIXEL_COUNT[3:0]]:
		({(VBORDER&HBORDER),(VBLANKING|HBLANKING)} == 2'b11)	?	BORDER[1]:
																					1'b0;

assign BLUE0X =	({VBLANKING,HBLANKING} == 2'b00)				?	BLUE0S[~PIXEL_COUNT[3:0]]:
		({(VBORDER&HBORDER),(VBLANKING|HBLANKING)} == 2'b11)	?	BORDER[0]:
																					1'b0;
/*****************************************************************************
* Switches to set different video modes
******************************************************************************/
assign MODE_256 = (COCO == 1'b1)					?	1'b1:
						({COCO, HRES[0]}== 2'b00)	?	1'b1:
																1'b0;

assign LINES_ROW	=	(~COCO)	?	LPR:
		({COCO, V} == 4'b1001)	?	3'b010:			// 3
		({COCO, V} == 4'b1010)	?	3'b010:			// 3
		({COCO, V} == 4'b1011)	?	3'b001:			// 2
		({COCO, V} == 4'b1100)	?	3'b001:			// 2
		({COCO, V} == 4'b1101)	?	3'b000:			// 1
		({COCO, V} == 4'b1110)	?	3'b000:			// 1
											3'b110;			// 12
/*****************************************************************************
* Count pixels across each line
* 32 and 40 character modes use double wide pixels
******************************************************************************/
always @ (posedge PIX_CLK or negedge RESET_N)
begin
	if(~RESET_N)
	begin
		PIXEL_COUNT <= 10'd000;
		HBLANKING <= 1'b1;
		HSYNC <= 1'b1;
		SYNC_FLAG <= 1'b0;
		HBORDER <= 1'b1;
		READMEM <= 1'b0;
	end
	else
	begin
		case (PIXEL_COUNT[2:0])
		3'b000:
		begin
	      READMEM <= 1'b0;
			CHAR_LATCH3 <= CHAR_LATCH;
			ATRIB_LATCH3 <= ATRIB_LATCH;
			if(VBANK==1'b0)
			begin
				CHAR_LATCH <= RAM_DATA[7:0];
				ATRIB_LATCH <= RAM_DATA[15:8];
			end
			else
			begin
				CHAR_LATCH <= RAM_DATA[23:16];
				ATRIB_LATCH <= RAM_DATA[31:24];
			end
		end
		3'b111:
		      READMEM <= 1'b1;
		default:
		      READMEM <= 1'b0;
		endcase

		case (PIXEL_COUNT)
		10'd013:				// First character read
		begin
			PIXEL_COUNT <= 10'd014;
			HBORDER <= 1'b1;
		end
		10'd015:				// Turn off horizontal blanking so first character can be displayed
		begin
			HBLANKING <= 1'b0;							// Turn off blanking
			HBORDER <= 1'b1;
			HSYNC <= 1'b1;									// Not H Sync
			PIXEL_COUNT  <= 10'd016;					// Next step
		end
		10'd527:											// 512 + 16 -1
		begin
			HBORDER <= 1'b1;
			HSYNC <= 1'b1;							// Not H Sync
			if(MODE_256)								// 512 mode
			begin
				HBLANKING <= 1'b1;					// Turn on blanking
				PIXEL_COUNT  <= 10'd592;			// 528 + 64 = 528 + 128 - 64
			end
			else											// 640 mode
			begin
				HBLANKING <= 1'b0;					// Leave blanking off
				PIXEL_COUNT  <= 10'd528;
			end
		end
		10'd655:											// 640 + 16 - 1
		begin
			HBLANKING <= 1'b1;						// Blanking on
			HBORDER <= 1'b1;
			HSYNC <= 1'b1;								// Not H Sync
			PIXEL_COUNT  <= 10'd656;
		end
		10'd657:											// 648 + 24 - 1
		begin
			HBLANKING <= 1'b1;
			HBORDER <= 1'b0;
			HSYNC <= 1'b1;
			PIXEL_COUNT <= 10'd658;
		end
		10'd671:											// 648 + 24 - 1
		begin
			HBLANKING <= 1'b1;
			HBORDER <= 1'b0;
			HSYNC <= 1'b0;								// Turn on Sync
			PIXEL_COUNT <= 10'd672;
		end
		10'd767:											// 672 + 104 - 1
		begin
			HBLANKING <= 1'b1;
			HSYNC <= 1'b1;								// SYNC OFF
			if(~MODE_256)									// 640 mode
				PIXEL_COUNT <= 10'd832;				// skip 64
			else
				PIXEL_COUNT <= 10'd768;
		end
		10'd799:
		begin
			PIXEL_COUNT <= 10'd800;
			HBORDER <= 1'b1;
		end
		10'd863:											// 864 - 1
		begin
			PIXEL_COUNT <= 10'd000;
			HSYNC <= 1'b1;
			SYNC_FLAG <= ~SYNC_FLAG;
		end
		default:
		begin
			PIXEL_COUNT <= PIXEL_COUNT + 1'b1;
		end
		endcase
	end
end

/*****************************************************************************
* Keeps track of how many rows are in each field.
******************************************************************************/
always @ (negedge ROW or posedge VBLANKING)
begin
	if(VBLANKING)
	begin
		VADD <= 8'h00;							// modify this to calculate the starting address
		if(COCO)
		begin
			ROW_ADD <= {SCRN_START_MSB[7:5],VERT,SCRN_START_LSB[5:0],3'h0};
		end
		else
		begin
			ROW_ADD <= {SCRN_START_MSB,SCRN_START_LSB,3'h0} + {HOR_OFFSET, 1'b0};
		end
	end
	else
	begin
		VADD <= VADD + 1'b1;					// modify this to add the line increment.
		ROW_ADD <= START_ADD;
	end
end

/*****************************************************************************
* Keeps track of how many lines are in each row.
* There are 2X lines per coco line.
******************************************************************************/
always @ (negedge HSYNC)
begin
	if(VBLANKING)
	begin
		if(~COCO)
			VLPR <= {VERT_FIN_SCRL, 1'b0};
		else
			VLPR <= 5'd0;
		ROW <= 1'b0;
		SIX <= 1'b0;
	end
	else
	begin
		case (VLPR)
		5'd0:										//Pixel Row 0
		begin
			VLPR <= 5'd01;
			if(LINES_ROW == 3'b000)			// 1
				ROW <= 1'b1;
			else
				ROW <= 1'b0;
		end
		5'd1:										//Pixel Row 0
		begin
			ROW <= 1'b0;
			if(LINES_ROW == 3'b000)			// 1
				VLPR <= 5'd0;
			else
				VLPR <= 5'd2;
		end
		5'd2:										//Pixel Row 1
		begin
			VLPR <= 5'd3;
			if(LINES_ROW == 3'b001)				// 2
				ROW <= 1'b1;
			else
				ROW <= 1'b0;
		end
		5'd3:										//Pixel Row 1
		begin
			ROW <= 1'b0;
			if(LINES_ROW == 3'b001)				// 2
				VLPR <= 5'd0;
			else
				VLPR <= 5'd4;
		end
		5'd4:										//Pixel Row 2
		begin
			VLPR <= 5'd5;
			if(LINES_ROW == 3'b010)				// 3
				ROW <= 1'b1;
			else
				ROW <= 1'b0;
		end
		5'd5:										//Pixel Row 2
		begin
			ROW <= 1'b0;
			if(LINES_ROW == 3'b010)				// 3
				VLPR <= 5'd0;
			else
				VLPR <= 5'd6;
		end
		5'd11:									//Pixel Row 5
		begin
			SIX <= 1'b1;
			VLPR <= 5'd12;
		end
		5'd13:									// Pixel Row 6
		begin
			VLPR <= 5'd14;
			if(LINES_ROW == 3'b011)			// 8
				ROW <= 1'b1;
			else
				ROW <= 1'b0;
		end
		5'd15:									// Pixel Row 7
		begin
			if(LINES_ROW == 3'b011)			// 8
			begin
				ROW <= 1'b0;
				SIX <= 1'b0;
				VLPR <= 5'd0;
			end
			else
			begin
				VLPR <= 5'd16;
				if(LINES_ROW == 3'b100)			// 9
					ROW <= 1'b1;
				else
					ROW <= 1'b0;
			end
		end
		5'd17:
		begin
			if(LINES_ROW == 3'b100)				// 9
			begin
				ROW <= 1'b0;
				SIX <= 1'b0;
				VLPR <= 5'd0;
			end
			else
			begin
				VLPR <= 5'd18;
				if(LINES_ROW == 3'b101)			// 10
					ROW <= 1'b1;
				else
					ROW <= 1'b0;
			end
		end
		5'd19:
		begin
			if(LINES_ROW == 3'b101)		// 10
			begin
				ROW <= 1'b0;
				VLPR <= 5'd0;
				SIX <= 1'b0;
			end
			else
				VLPR <= 5'd20;
		end
		5'd21:
		begin
			VLPR <= 5'd22;
			if(LINES_ROW == 3'b110)				// 12
				ROW <= 1'b1;
			else
				ROW <= 1'b0;
		end
		5'd23:						// 12 *2 -1 = 23 = 0x17
		begin
			ROW <= 1'b0;
			SIX <= 1'b0;
			if(LINES_ROW == 3'b110)		// 12
				VLPR <= 5'd0;
			else
				VLPR <= 5'd24;
		end
//		5'd30:						// 12 *2 -1 = 23 = 0x17
//		begin
//			ROW <= 1'b1;
//			VLPR <= 5'd31;
//		end
		5'd31:						// 16 *2 -1 = 31 = 0x1F
		begin
			if(LINES_ROW == 3'b111)				// 1/0
				VLPR <= 5'd31;
			else
			begin
				VLPR <= 5'd0;
			end
		end
		default:
			VLPR <= VLPR + 1'b1;
		endcase
	end
end

/*****************************************************************************
* Keeps track of the real line number, and controls VSYNC and VBlanking.
* Does not keep track of the lines per row
*
*	LPR				Lines
*
*	00 or COCO =1	192
*	01					200
*	10					210
*	11					225	(25*9)
******************************************************************************/
always @ (negedge HSYNC or negedge RESET_N)
begin
	if(~RESET_N)
	begin
		LINE <= 10'd00;
		VBLANKING <= 1'b0;
		VSYNC <= 1'b1;
	end
	else
	case (LINE)
	10'd383:								// End of 192 line display
	begin
		LINE <= 10'd384;
		VSYNC <= 1'b1;
		VBORDER <= 1'b1;
		if((LPF == 2'b00) || (COCO == 1'b1))		// Standard COCO modes are always 192
		begin
			VBLANKING <= 1'b1;
		end
	end
	10'd399:								// End of 200 line display
	begin
		LINE <= 10'd400;
		VSYNC <= 1'b1;
		VBORDER <= 1'b1;
		if(LPF == 2'b01)
		begin
			VBLANKING <= 1'b1;
		end
	end
	10'd419:								// End of 210 line display
	begin
		LINE <= 10'd420;
		VSYNC <= 1'b1;
		VBORDER <= 1'b1;
		if(LPF == 2'b10)
		begin
			VBLANKING <= 1'b1;
		end
	end
	10'd449:								// End of 225 line display
	begin
		LINE <= 10'd450;
		VSYNC <= 1'b1;
		VBLANKING <= 1'b1;
		VBORDER <= 1'b1;
	end
	10'd457:
	begin
		VBORDER <= 1'b0;
		LINE <= 10'd458;
	end
// 10'd432:	Start Clock
// 10'd439:	Stop Clock and end border color
	10'd469:
	begin
		LINE <= 10'd470;
		VSYNC <= 1'b0;					// Sync on
		VBLANKING <= 1'b1;
		VBORDER <= 1'b0;
	end
	10'd471:
	begin
		LINE <= 10'd472;
		VSYNC <= 1'b1;					// Sync off
		VBLANKING <= 1'b1;
		VBORDER <= 1'b0;
	end
	10'd512:
	begin
		LINE <= 10'd513;
		VBLANKING <= 1'b1;
		VBORDER <= 1'b1;
		VSYNC <= 1'b1;
	end
	10'd520:							// -1
	begin
		LINE <= 10'd000;
		VBLANKING <= 1'b0;
		VBORDER <= 1'b1;
		VSYNC <= 1'b1;
	end
	default:
	begin
		LINE <= LINE + 1'b1;
	end
	endcase
end
endmodule
