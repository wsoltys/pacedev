library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.project_pkg.all;
use work.target_pkg.all;

package platform_pkg is

	--  
	-- PACE constants which *MUST* be defined
	--
	
	constant PACE_VIDEO_NUM_BITMAPS		    : natural := 0;
	constant PACE_VIDEO_NUM_TILEMAPS	    : natural := 1;
	constant PACE_VIDEO_NUM_SPRITES 	    : natural := 0;
	constant PACE_VIDEO_H_SIZE				    : integer := 256;
	constant PACE_VIDEO_V_SIZE				    : integer := 256;
  constant PACE_VIDEO_PIPELINE_DELAY    : integer := 5;
	
	constant PACE_INPUTS_NUM_BYTES        : integer := 3;
	
	--
	-- Platform-specific constants (optional)
	--

	constant CABAL_1MHz_CLK0_COUNTS			    : natural := 
    PACE_CLKIN0 * PACE_CLK0_MULTIPLY_BY / PACE_CLK0_DIVIDE_BY;

	constant CABAL_CPU_CLK_ENA_DIVIDE_BY	  : natural := 
    CABAL_1MHz_CLK0_COUNTS / 3;

  constant CABAL_SRC_DIR                  : string;

	-- Palette : Table of RGB entries	

	type pal_entry_typ is array (0 to 2) of std_logic_vector(5 downto 0);
	type pal_typ is array (0 to 255) of pal_entry_typ;

	constant pal : pal_typ :=
	(
		0 => (0=>"111100", 1=>"101111", 2=>"100011"),
		1 => (0=>"111000", 1=>"100011", 2=>"000000"),
		2 => (0=>"110100", 1=>"000000", 2=>"000000"),
		4 => (0=>"111111", 1=>"111111", 2=>"111111"),
		5 => (0=>"000000", 1=>"000000", 2=>"111111"),
		6 => (0=>"111111", 1=>"000000", 2=>"000000"),
		8 => (0=>"000000", 1=>"000000", 2=>"111000"),
		9 => (0=>"101111", 1=>"010100", 2=>"000000"),
		10 => (0=>"111000", 1=>"000000", 2=>"000000"),
		12 => (0=>"111111", 1=>"000000", 2=>"000000"),
		13 => (0=>"000000", 1=>"000000", 2=>"111111"),
		14 => (0=>"000000", 1=>"100111", 2=>"000000"),
		16 => (0=>"111111", 1=>"111111", 2=>"111111"),
		17 => (0=>"000000", 1=>"000000", 2=>"111111"),
		18 => (0=>"000000", 1=>"000000", 2=>"100111"),
		21 => (0=>"011100", 1=>"011100", 2=>"011100"),
		22 => (0=>"100111", 1=>"100111", 2=>"100111"),
		24 => (0=>"111111", 1=>"111111", 2=>"111111"),
		25 => (0=>"111111", 1=>"111111", 2=>"111111"),
		26 => (0=>"110100", 1=>"011000", 2=>"001011"),
		28 => (0=>"000000", 1=>"011100", 2=>"101111"),
		29 => (0=>"000000", 1=>"011100", 2=>"101111"),
		30 => (0=>"000000", 1=>"101111", 2=>"111000"),
		32 => (0=>"111000", 1=>"000000", 2=>"010100"),
		33 => (0=>"111000", 1=>"000000", 2=>"010100"),
		34 => (0=>"111111", 1=>"110100", 2=>"010000"),
		37 => (0=>"110100", 1=>"111100", 2=>"111111"),
		38 => (0=>"101111", 1=>"110100", 2=>"111100"),
		40 => (0=>"111100", 1=>"000000", 2=>"000000"),
		41 => (0=>"000000", 1=>"000000", 2=>"100011"),
		42 => (0=>"000000", 1=>"000000", 2=>"111100"),
		68 => (0=>"000011", 1=>"000011", 2=>"000011"),
		72 => (0=>"000111", 1=>"000111", 2=>"000111"),
		76 => (0=>"001011", 1=>"001011", 2=>"001011"),
		80 => (0=>"010000", 1=>"010000", 2=>"010000"),
		84 => (0=>"010100", 1=>"010100", 2=>"010100"),
		88 => (0=>"011000", 1=>"011000", 2=>"011000"),
		92 => (0=>"011100", 1=>"011100", 2=>"011100"),
		96 => (0=>"100011", 1=>"100011", 2=>"100011"),
		100 => (0=>"100111", 1=>"100111", 2=>"100111"),
		104 => (0=>"101011", 1=>"101011", 2=>"101011"),
		108 => (0=>"101111", 1=>"101111", 2=>"101111"),
		112 => (0=>"110100", 1=>"110100", 2=>"110100"),
		116 => (0=>"111000", 1=>"111000", 2=>"111000"),
		120 => (0=>"111100", 1=>"111100", 2=>"111100"),
		124 => (0=>"111111", 1=>"111111", 2=>"111111"),
		128 => (0=>"000000", 1=>"001011", 2=>"011000"),
		129 => (0=>"111111", 1=>"111000", 2=>"011100"),
		130 => (0=>"110100", 1=>"101011", 2=>"000000"),
		132 => (0=>"000000", 1=>"001011", 2=>"011000"),
		133 => (0=>"111111", 1=>"111111", 2=>"111111"),
		134 => (0=>"111000", 1=>"000000", 2=>"000000"),
		136 => (0=>"000000", 1=>"001011", 2=>"011000"),
		137 => (0=>"111111", 1=>"111000", 2=>"011100"),
		138 => (0=>"000000", 1=>"100111", 2=>"000000"),
		140 => (0=>"000000", 1=>"001011", 2=>"011000"),
		141 => (0=>"111111", 1=>"111111", 2=>"111111"),
		142 => (0=>"000000", 1=>"100111", 2=>"000000"),
		144 => (0=>"000000", 1=>"001011", 2=>"011000"),
		145 => (0=>"111111", 1=>"111000", 2=>"011100"),
		others => (others => (others => '0'))
	);

end;
