library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.project_pkg.all;
use work.target_pkg.all;
use work.platform_variant_pkg.all;

package platform_pkg is

	--  
	-- PACE constants which *MUST* be defined
	--

	constant PACE_VIDEO_NUM_BITMAPS		    : natural := 0;
	constant PACE_VIDEO_NUM_TILEMAPS 	    : natural := 2;
	constant PACE_VIDEO_NUM_SPRITES 	    : natural := 0;
	constant PACE_VIDEO_H_SIZE				    : integer := 256; -- clipped to 224
	constant PACE_VIDEO_V_SIZE				    : integer := 288;
  constant PACE_VIDEO_PIPELINE_DELAY    : integer := 3;
	
  constant PACE_INPUTS_NUM_BYTES        : integer := 3;

	constant CLK0_FREQ_MHz		            : natural := 
    PACE_CLKIN0 * PACE_CLK0_MULTIPLY_BY / PACE_CLK0_DIVIDE_BY;
  
	--
	-- Platform-specific constants (optional)
	--

  constant GALAGA_SOURCE_ROOT_DIR       : string := "../../../../../src/platform/galaga/";
  constant VARIANT_SOURCE_ROOT_DIR      : string := GALAGA_SOURCE_ROOT_DIR & 
                                                    PLATFORM_VARIANT & "/";
  constant VARIANT_ROM_DIR              : string := VARIANT_SOURCE_ROOT_DIR & 
                                                    "roms/";
  
	type pal_entry_typ is array (0 to 2) of std_logic_vector(5 downto 0);
	type pal_typ is array (0 to 127) of pal_entry_typ;

	constant pal : pal_typ :=
	(
    1 => (0=>"011000", 1=>"011000", 2=>"011000"),
    2 => (0=>"001011", 1=>"100011", 2=>"111111"),
    3 => (0=>"000000", 1=>"110100", 2=>"110100"),
    4 => (0=>"010100", 1=>"000111", 2=>"000111"),
    5 => (0=>"101011", 1=>"101011", 2=>"101011"),
    6 => (0=>"000111", 1=>"011100", 2=>"111111"),
    7 => (0=>"010100", 1=>"010000", 2=>"111111"),
    8 => (0=>"100111", 1=>"100111", 2=>"000000"),
    9 => (0=>"110100", 1=>"110100", 2=>"110100"),
    10 => (0=>"010000", 1=>"100011", 2=>"000111"),
    11 => (0=>"010000", 1=>"011000", 2=>"000000"),
    12 => (0=>"100111", 1=>"100111", 2=>"010000"),
    13 => (0=>"011000", 1=>"001011", 2=>"000111"),
    14 => (0=>"010100", 1=>"010100", 2=>"000111"),
    15 => (0=>"010100", 1=>"010100", 2=>"010100"),
    16 => (0=>"011100", 1=>"100011", 2=>"001011"),
    17 => (0=>"010100", 1=>"100011", 2=>"001011"),
    18 => (0=>"010100", 1=>"100011", 2=>"100111"),
    19 => (0=>"100011", 1=>"011000", 2=>"000000"),
    20 => (0=>"111000", 1=>"101111", 2=>"000000"),
    21 => (0=>"110100", 1=>"011000", 2=>"000000"),
    22 => (0=>"011100", 1=>"010000", 2=>"000000"),
    23 => (0=>"010000", 1=>"001011", 2=>"000111"),
    24 => (0=>"000111", 1=>"000111", 2=>"000000"),
    25 => (0=>"000111", 1=>"010000", 2=>"000000"),
    26 => (0=>"000111", 1=>"011000", 2=>"000000"),
    27 => (0=>"001011", 1=>"011100", 2=>"000011"),
    28 => (0=>"010100", 1=>"100111", 2=>"110100"),
    29 => (0=>"100111", 1=>"100111", 2=>"011100"),
    30 => (0=>"011100", 1=>"100011", 2=>"000111"),
    31 => (0=>"100011", 1=>"100011", 2=>"000111"),
    32 => (0=>"101011", 1=>"100011", 2=>"010000"),
    33 => (0=>"100011", 1=>"011000", 2=>"000111"),
    34 => (0=>"011100", 1=>"011000", 2=>"000000"),
    35 => (0=>"011000", 1=>"010100", 2=>"000000"),
    36 => (0=>"011100", 1=>"011100", 2=>"011100"),
    37 => (0=>"100011", 1=>"100011", 2=>"100011"),
    38 => (0=>"111111", 1=>"000000", 2=>"000000"),
    39 => (0=>"010000", 1=>"100011", 2=>"011100"),
    40 => (0=>"001011", 1=>"011100", 2=>"101111"),
    41 => (0=>"000000", 1=>"100011", 2=>"110100"),
    42 => (0=>"111000", 1=>"101111", 2=>"011000"),
    43 => (0=>"000000", 1=>"011000", 2=>"100011"),
    44 => (0=>"101011", 1=>"101111", 2=>"110100"),
    45 => (0=>"000111", 1=>"010100", 2=>"101011"),
    46 => (0=>"000000", 1=>"110100", 2=>"000000"),
    47 => (0=>"101011", 1=>"000000", 2=>"000000"),
    48 => (0=>"000111", 1=>"010000", 2=>"011000"),
    49 => (0=>"010000", 1=>"100011", 2=>"101111"),
    50 => (0=>"010100", 1=>"010100", 2=>"000000"),
    51 => (0=>"101011", 1=>"101011", 2=>"000000"),
    52 => (0=>"100011", 1=>"100011", 2=>"011000"),
    53 => (0=>"100011", 1=>"010000", 2=>"010000"),
    54 => (0=>"111111", 1=>"111111", 2=>"000000"),
    55 => (0=>"111111", 1=>"101011", 2=>"000000"),
    56 => (0=>"111111", 1=>"011000", 2=>"000000"),
    57 => (0=>"000111", 1=>"011000", 2=>"101011"),
    58 => (0=>"111100", 1=>"101011", 2=>"000000"),
    59 => (0=>"110100", 1=>"000000", 2=>"000000"),
    60 => (0=>"000000", 1=>"000000", 2=>"111111"),
    61 => (0=>"111111", 1=>"111111", 2=>"111111"),
    62 => (0=>"111100", 1=>"111100", 2=>"111100"),
    63 => (0=>"000111", 1=>"000111", 2=>"000111"),
    64 => (0=>"110100", 1=>"011000", 2=>"000000"),
    65 => (0=>"111000", 1=>"101111", 2=>"000000"),
    66 => (0=>"000000", 1=>"010100", 2=>"000000"),
    67 => (0=>"000000", 1=>"100011", 2=>"000000"),
    68 => (0=>"010000", 1=>"010000", 2=>"010000"),
    69 => (0=>"000000", 1=>"111111", 2=>"111111"),
    70 => (0=>"000000", 1=>"100011", 2=>"111111"),
    71 => (0=>"100011", 1=>"000000", 2=>"000000"),
    72 => (0=>"011000", 1=>"000000", 2=>"000000"),
    73 => (0=>"000000", 1=>"001011", 2=>"000000"),
    74 => (0=>"110100", 1=>"010000", 2=>"011000"),
    75 => (0=>"010000", 1=>"010000", 2=>"011000"),
    76 => (0=>"010100", 1=>"010100", 2=>"100011"),
    77 => (0=>"100011", 1=>"100011", 2=>"101011"),
    78 => (0=>"011100", 1=>"011100", 2=>"100111"),
    79 => (0=>"011000", 1=>"011000", 2=>"100011"),
    80 => (0=>"000111", 1=>"000111", 2=>"100011"),
    81 => (0=>"100011", 1=>"011000", 2=>"000111"),
    82 => (0=>"000111", 1=>"010100", 2=>"101111"),
    83 => (0=>"010100", 1=>"010000", 2=>"000000"),
    84 => (0=>"101111", 1=>"011100", 2=>"000111"),
    85 => (0=>"111111", 1=>"100011", 2=>"111111"),
    86 => (0=>"110100", 1=>"010000", 2=>"010000"),
    87 => (0=>"000000", 1=>"110100", 2=>"111111"),
    88 => (0=>"101011", 1=>"011000", 2=>"000000"),
    89 => (0=>"010000", 1=>"000000", 2=>"000000"),
    90 => (0=>"111100", 1=>"111100", 2=>"000000"),
    91 => (0=>"111111", 1=>"110100", 2=>"101011"),
    92 => (0=>"111111", 1=>"110100", 2=>"011000"),
    93 => (0=>"111111", 1=>"110100", 2=>"010000"),
    94 => (0=>"110100", 1=>"100011", 2=>"010000"),
    95 => (0=>"110100", 1=>"110100", 2=>"110100"),
    96 => (0=>"111111", 1=>"111111", 2=>"011000"),
    97 => (0=>"101111", 1=>"101111", 2=>"010000"),
    98 => (0=>"011100", 1=>"011100", 2=>"000111"),
    99 => (0=>"001011", 1=>"001011", 2=>"001011"),
    100 => (0=>"111111", 1=>"100011", 2=>"000000"),
    101 => (0=>"010000", 1=>"010000", 2=>"110100"),
    102 => (0=>"010000", 1=>"010000", 2=>"000111"),
    103 => (0=>"011000", 1=>"011000", 2=>"010000"),
    104 => (0=>"101011", 1=>"101011", 2=>"100011"),
    105 => (0=>"110100", 1=>"110100", 2=>"101011"),
    106 => (0=>"101011", 1=>"100011", 2=>"010000"),
    107 => (0=>"100011", 1=>"010000", 2=>"000111"),
    108 => (0=>"000000", 1=>"111111", 2=>"000000"),
    109 => (0=>"100011", 1=>"000000", 2=>"111111"),
    110 => (0=>"111111", 1=>"000000", 2=>"111111"),
    111 => (0=>"100011", 1=>"010000", 2=>"000000"),
    112 => (0=>"010000", 1=>"000111", 2=>"000000"),
    113 => (0=>"100011", 1=>"100011", 2=>"000000"),
    114 => (0=>"010000", 1=>"010000", 2=>"000000"),
    115 => (0=>"000000", 1=>"010000", 2=>"000000"),
    116 => (0=>"000000", 1=>"100011", 2=>"100011"),
    117 => (0=>"000000", 1=>"010000", 2=>"010000"),
    118 => (0=>"000000", 1=>"000000", 2=>"100011"),
    119 => (0=>"000000", 1=>"000000", 2=>"010000"),
    120 => (0=>"010000", 1=>"000000", 2=>"100011"),
    121 => (0=>"000111", 1=>"000000", 2=>"010000"),
    122 => (0=>"100011", 1=>"000000", 2=>"100011"),
    123 => (0=>"010000", 1=>"000000", 2=>"010000"),
    124 => (0=>"111111", 1=>"111111", 2=>"110100"),
    125 => (0=>"111111", 1=>"111111", 2=>"101011"),
    126 => (0=>"111111", 1=>"101011", 2=>"011000"),
		others => (others => (others => '0'))
	);

	-- Colour Look-up Table (CLUT) : Table of palette entries
	-- - each row has four (4) palette indexes
	--   decoded from 2 bits of tile data
	
	type clut_entry_typ is array (0 to 3) of std_logic_vector(3 downto 0);
	type clut_typ is array (0 to 63) of clut_entry_typ;

	constant clut : clut_typ :=
	(
		1 => (0=>X"0", 1=>X"5", 2=>X"3", 3=>X"1"),
		2 => (0=>X"0", 1=>X"5", 2=>X"2", 3=>X"1"),
		3 => (0=>X"0", 1=>X"5", 2=>X"6", 3=>X"1"),
		4 => (0=>X"0", 1=>X"5", 2=>X"7", 3=>X"1"),
		5 => (0=>X"0", 1=>X"5", 2=>X"A", 3=>X"1"),
		6 => (0=>X"0", 1=>X"5", 2=>X"B", 3=>X"1"),
		7 => (0=>X"0", 1=>X"5", 2=>X"C", 3=>X"1"),
		8 => (0=>X"0", 1=>X"5", 2=>X"D", 3=>X"1"),
		9 => (0=>X"0", 1=>X"5", 2=>X"4", 3=>X"1"),
		10 => (0=>X"0", 1=>X"3", 2=>X"6", 3=>X"1"),
		11 => (0=>X"0", 1=>X"3", 2=>X"2", 3=>X"1"),
		12 => (0=>X"0", 1=>X"3", 2=>X"7", 3=>X"1"),
		13 => (0=>X"0", 1=>X"3", 2=>X"5", 3=>X"1"),
		14 => (0=>X"0", 1=>X"2", 2=>X"3", 3=>X"1"),
		16 => (0=>X"0", 1=>X"8", 2=>X"3", 3=>X"1"),
		17 => (0=>X"0", 1=>X"9", 2=>X"2", 3=>X"5"),
		18 => (0=>X"0", 1=>X"8", 2=>X"5", 3=>X"D"),
		19 => (0=>X"4", 1=>X"4", 2=>X"4", 3=>X"4"),
		22 => (0=>X"0", 1=>X"2", 2=>X"2", 3=>X"2"),
		23 => (0=>X"0", 1=>X"3", 2=>X"3", 3=>X"3"),
		24 => (0=>X"0", 1=>X"6", 2=>X"6", 3=>X"6"),
		25 => (0=>X"0", 1=>X"7", 2=>X"7", 3=>X"7"),
		26 => (0=>X"0", 1=>X"A", 2=>X"A", 3=>X"A"),
		27 => (0=>X"0", 1=>X"B", 2=>X"B", 3=>X"B"),
		28 => (0=>X"0", 1=>X"1", 2=>X"1", 3=>X"1"),
		29 => (0=>X"0", 1=>X"5", 2=>X"5", 3=>X"5"),
		30 => (0=>X"8", 1=>X"9", 2=>X"A", 3=>X"B"),
		31 => (0=>X"C", 1=>X"D", 2=>X"E", 3=>X"F"),
		33 => (0=>X"0", 1=>X"3", 2=>X"7", 3=>X"D"),
		34 => (0=>X"0", 1=>X"C", 2=>X"F", 3=>X"B"),
		35 => (0=>X"0", 1=>X"C", 2=>X"E", 3=>X"B"),
		36 => (0=>X"0", 1=>X"C", 2=>X"6", 3=>X"B"),
		37 => (0=>X"0", 1=>X"C", 2=>X"7", 3=>X"B"),
		38 => (0=>X"0", 1=>X"C", 2=>X"3", 3=>X"B"),
		39 => (0=>X"0", 1=>X"C", 2=>X"8", 3=>X"B"),
		40 => (0=>X"0", 1=>X"C", 2=>X"D", 3=>X"B"),
		41 => (0=>X"0", 1=>X"C", 2=>X"4", 3=>X"B"),
		42 => (0=>X"0", 1=>X"C", 2=>X"9", 3=>X"B"),
		43 => (0=>X"0", 1=>X"C", 2=>X"5", 3=>X"B"),
		44 => (0=>X"0", 1=>X"C", 2=>X"2", 3=>X"B"),
		45 => (0=>X"0", 1=>X"C", 2=>X"B", 3=>X"2"),
		46 => (0=>X"0", 1=>X"8", 2=>X"C", 3=>X"2"),
		47 => (0=>X"0", 1=>X"8", 2=>X"F", 3=>X"2"),
		48 => (0=>X"0", 1=>X"3", 2=>X"2", 3=>X"1"),
		49 => (0=>X"0", 1=>X"2", 2=>X"F", 3=>X"3"),
		50 => (0=>X"0", 1=>X"F", 2=>X"E", 3=>X"2"),
		51 => (0=>X"0", 1=>X"E", 2=>X"7", 3=>X"F"),
		52 => (0=>X"0", 1=>X"7", 2=>X"6", 3=>X"E"),
		53 => (0=>X"0", 1=>X"6", 2=>X"5", 3=>X"7"),
		54 => (0=>X"0", 1=>X"5", 2=>X"0", 3=>X"6"),
		55 => (0=>X"0", 1=>X"0", 2=>X"B", 3=>X"5"),
		56 => (0=>X"0", 1=>X"B", 2=>X"C", 3=>X"0"),
		57 => (0=>X"0", 1=>X"C", 2=>X"D", 3=>X"B"),
		58 => (0=>X"0", 1=>X"D", 2=>X"8", 3=>X"C"),
		59 => (0=>X"0", 1=>X"8", 2=>X"9", 3=>X"D"),
		60 => (0=>X"0", 1=>X"9", 2=>X"A", 3=>X"8"),
		61 => (0=>X"0", 1=>X"A", 2=>X"1", 3=>X"9"),
		62 => (0=>X"0", 1=>X"1", 2=>X"4", 3=>X"A"),
		63 => (0=>X"0", 1=>X"4", 2=>X"3", 3=>X"1"),
		others => (others => (others => '0'))
	);


  type from_PLATFORM_IO_t is record
    not_used  : std_logic;
  end record;

  type to_PLATFORM_IO_t is record
    not_used  : std_logic;
  end record;

end;
