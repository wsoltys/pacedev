library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

package platform_variant_pkg is

	--
	-- Platform-variant-specific constants (optional)
	--

  constant PLATFORM_VARIANT         : string := "mac128k";
  
end;
