-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_PGM_67 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_PGM_67 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"6F",x"7E",x"2C",x"66",x"6F",x"22",x"82",x"83", -- 0x0000
    x"18",x"13",x"32",x"2F",x"84",x"CD",x"F9",x"07", -- 0x0008
    x"21",x"40",x"B0",x"01",x"00",x"18",x"71",x"2C", -- 0x0010
    x"10",x"FC",x"CD",x"45",x"38",x"3E",x"20",x"32", -- 0x0018
    x"6A",x"82",x"3E",x"80",x"DF",x"21",x"44",x"80", -- 0x0020
    x"AF",x"77",x"23",x"77",x"23",x"77",x"23",x"36", -- 0x0028
    x"F0",x"D1",x"E1",x"AF",x"32",x"9B",x"82",x"32", -- 0x0030
    x"EA",x"83",x"32",x"4D",x"82",x"32",x"49",x"82", -- 0x0038
    x"32",x"51",x"82",x"3C",x"32",x"6C",x"82",x"32", -- 0x0040
    x"CD",x"83",x"3E",x"10",x"32",x"68",x"82",x"C9", -- 0x0048
    x"3A",x"6C",x"82",x"A7",x"C8",x"21",x"6A",x"82", -- 0x0050
    x"35",x"C0",x"AF",x"32",x"6C",x"82",x"C9",x"3A", -- 0x0058
    x"47",x"80",x"FE",x"30",x"D8",x"FE",x"D0",x"4F", -- 0x0060
    x"28",x"17",x"D0",x"3A",x"69",x"82",x"B9",x"D8", -- 0x0068
    x"C8",x"79",x"32",x"69",x"82",x"11",x"01",x"00", -- 0x0070
    x"FE",x"80",x"C8",x"E5",x"CD",x"03",x"09",x"E1", -- 0x0078
    x"C9",x"3A",x"69",x"82",x"A7",x"20",x"E4",x"3E", -- 0x0080
    x"E0",x"32",x"69",x"82",x"18",x"DD",x"DD",x"21", -- 0x0088
    x"73",x"82",x"DD",x"7E",x"02",x"32",x"1A",x"81", -- 0x0090
    x"3A",x"10",x"81",x"3C",x"32",x"10",x"81",x"FE", -- 0x0098
    x"50",x"D4",x"84",x"31",x"DD",x"21",x"7C",x"82", -- 0x00A0
    x"DD",x"7E",x"02",x"32",x"19",x"81",x"3A",x"11", -- 0x00A8
    x"81",x"3C",x"3C",x"32",x"11",x"81",x"FE",x"A0", -- 0x00B0
    x"DC",x"25",x"32",x"3A",x"6E",x"82",x"3C",x"32", -- 0x00B8
    x"6E",x"82",x"FE",x"10",x"CA",x"D2",x"30",x"FE", -- 0x00C0
    x"20",x"CA",x"F8",x"30",x"FE",x"30",x"CA",x"1E", -- 0x00C8
    x"31",x"C9",x"21",x"73",x"82",x"7E",x"23",x"46", -- 0x00D0
    x"21",x"1A",x"81",x"4E",x"11",x"AC",x"24",x"32", -- 0x00D8
    x"B1",x"81",x"CD",x"55",x"31",x"21",x"7C",x"82", -- 0x00E0
    x"7E",x"23",x"46",x"21",x"19",x"81",x"4E",x"11", -- 0x00E8
    x"E8",x"24",x"32",x"B1",x"81",x"C3",x"48",x"31", -- 0x00F0
    x"21",x"73",x"82",x"7E",x"23",x"46",x"21",x"1A", -- 0x00F8
    x"81",x"4E",x"11",x"B4",x"24",x"32",x"B1",x"81", -- 0x0100
    x"CD",x"55",x"31",x"21",x"7C",x"82",x"7E",x"23", -- 0x0108
    x"46",x"21",x"19",x"81",x"4E",x"11",x"FC",x"24", -- 0x0110
    x"32",x"B1",x"81",x"C3",x"48",x"31",x"21",x"73", -- 0x0118
    x"82",x"7E",x"23",x"46",x"21",x"1A",x"81",x"4E", -- 0x0120
    x"11",x"BC",x"24",x"32",x"B1",x"81",x"AF",x"32", -- 0x0128
    x"6E",x"82",x"CD",x"55",x"31",x"21",x"7C",x"82", -- 0x0130
    x"7E",x"23",x"46",x"21",x"19",x"81",x"4E",x"11", -- 0x0138
    x"10",x"25",x"32",x"B1",x"81",x"C3",x"48",x"31", -- 0x0140
    x"2A",x"7E",x"24",x"ED",x"53",x"01",x"80",x"78", -- 0x0148
    x"32",x"03",x"80",x"18",x"0B",x"2A",x"78",x"24", -- 0x0150
    x"ED",x"53",x"01",x"80",x"78",x"32",x"03",x"80", -- 0x0158
    x"1A",x"77",x"23",x"13",x"1A",x"77",x"2B",x"D5", -- 0x0160
    x"11",x"20",x"00",x"19",x"D1",x"13",x"10",x"F0", -- 0x0168
    x"3A",x"B1",x"81",x"5F",x"16",x"00",x"19",x"3A", -- 0x0170
    x"03",x"80",x"47",x"ED",x"5B",x"01",x"80",x"0D", -- 0x0178
    x"C2",x"60",x"31",x"C9",x"DD",x"21",x"73",x"82", -- 0x0180
    x"AF",x"67",x"DD",x"46",x"01",x"C6",x"20",x"10", -- 0x0188
    x"FC",x"4F",x"DD",x"6E",x"00",x"09",x"5D",x"54", -- 0x0190
    x"AF",x"6F",x"67",x"DD",x"46",x"02",x"05",x"19", -- 0x0198
    x"10",x"FD",x"11",x"08",x"A8",x"19",x"0E",x"02", -- 0x01A0
    x"3A",x"10",x"81",x"FE",x"50",x"CA",x"C7",x"31", -- 0x01A8
    x"FE",x"80",x"CA",x"D5",x"31",x"FE",x"A0",x"CA", -- 0x01B0
    x"EE",x"31",x"FE",x"B0",x"CA",x"D5",x"31",x"FE", -- 0x01B8
    x"D0",x"CA",x"C7",x"31",x"C3",x"11",x"32",x"06", -- 0x01C0
    x"02",x"11",x"19",x"32",x"CD",x"01",x"32",x"0D", -- 0x01C8
    x"20",x"F5",x"C3",x"11",x"32",x"06",x"02",x"11", -- 0x01D0
    x"1D",x"32",x"CD",x"01",x"32",x"0D",x"20",x"F5", -- 0x01D8
    x"3A",x"07",x"81",x"A7",x"CA",x"11",x"32",x"AF", -- 0x01E0
    x"32",x"07",x"81",x"C3",x"11",x"32",x"06",x"02", -- 0x01E8
    x"11",x"21",x"32",x"CD",x"01",x"32",x"0D",x"20", -- 0x01F0
    x"F5",x"3E",x"01",x"32",x"07",x"81",x"C3",x"11", -- 0x01F8
    x"32",x"1A",x"77",x"13",x"23",x"1A",x"77",x"13", -- 0x0200
    x"D5",x"11",x"1F",x"00",x"19",x"D1",x"10",x"F1", -- 0x0208
    x"C9",x"DD",x"7E",x"02",x"3D",x"32",x"1A",x"81", -- 0x0210
    x"C9",x"94",x"95",x"96",x"97",x"98",x"99",x"9A", -- 0x0218
    x"9B",x"10",x"10",x"10",x"10",x"DD",x"21",x"7C", -- 0x0220
    x"82",x"AF",x"67",x"DD",x"46",x"01",x"C6",x"20", -- 0x0228
    x"10",x"FC",x"4F",x"DD",x"6E",x"00",x"09",x"5D", -- 0x0230
    x"54",x"AF",x"6F",x"67",x"DD",x"46",x"02",x"05", -- 0x0238
    x"19",x"10",x"FD",x"11",x"0E",x"A8",x"19",x"0E", -- 0x0240
    x"03",x"3A",x"11",x"81",x"FE",x"00",x"CA",x"68", -- 0x0248
    x"32",x"FE",x"30",x"CA",x"76",x"32",x"FE",x"50", -- 0x0250
    x"CA",x"8F",x"32",x"FE",x"60",x"CA",x"76",x"32", -- 0x0258
    x"FE",x"70",x"CA",x"68",x"32",x"C3",x"B2",x"32", -- 0x0260
    x"06",x"02",x"11",x"BA",x"32",x"CD",x"A2",x"32", -- 0x0268
    x"0D",x"20",x"F5",x"C3",x"B2",x"32",x"06",x"02", -- 0x0270
    x"11",x"BE",x"32",x"CD",x"A2",x"32",x"0D",x"20", -- 0x0278
    x"F5",x"3A",x"08",x"81",x"A7",x"CA",x"B2",x"32", -- 0x0280
    x"AF",x"32",x"08",x"81",x"C3",x"B2",x"32",x"06", -- 0x0288
    x"02",x"11",x"C2",x"32",x"CD",x"A2",x"32",x"0D", -- 0x0290
    x"20",x"F5",x"3E",x"01",x"32",x"08",x"81",x"C3", -- 0x0298
    x"B2",x"32",x"1A",x"77",x"13",x"23",x"1A",x"77", -- 0x02A0
    x"13",x"D5",x"11",x"1F",x"00",x"19",x"D1",x"10", -- 0x02A8
    x"F1",x"C9",x"DD",x"7E",x"02",x"3D",x"32",x"19", -- 0x02B0
    x"81",x"C9",x"94",x"95",x"96",x"97",x"98",x"99", -- 0x02B8
    x"9A",x"9B",x"10",x"10",x"10",x"10",x"D9",x"21", -- 0x02C0
    x"93",x"82",x"3A",x"FD",x"83",x"3D",x"28",x"01", -- 0x02C8
    x"2C",x"7E",x"01",x"E9",x"32",x"26",x"00",x"6F", -- 0x02D0
    x"85",x"6F",x"09",x"5E",x"23",x"56",x"EB",x"11", -- 0x02D8
    x"70",x"82",x"01",x"21",x"00",x"ED",x"B0",x"D9", -- 0x02E0
    x"C9",x"F3",x"32",x"14",x"33",x"35",x"33",x"56", -- 0x02E8
    x"33",x"77",x"33",x"60",x"08",x"03",x"60",x"04", -- 0x02F0
    x"04",x"80",x"0C",x"02",x"80",x"06",x"03",x"40", -- 0x02F8
    x"06",x"04",x"80",x"02",x"04",x"E0",x"04",x"02", -- 0x0300
    x"60",x"02",x"01",x"C0",x"02",x"03",x"C0",x"02", -- 0x0308
    x"03",x"E0",x"02",x"03",x"60",x"08",x"03",x"40", -- 0x0310
    x"04",x"05",x"80",x"0C",x"01",x"60",x"06",x"03", -- 0x0318
    x"C0",x"06",x"03",x"80",x"02",x"04",x"E0",x"04", -- 0x0320
    x"03",x"60",x"02",x"02",x"E0",x"02",x"04",x"C0", -- 0x0328
    x"02",x"04",x"E0",x"02",x"04",x"60",x"08",x"02", -- 0x0330
    x"80",x"04",x"04",x"80",x"0C",x"01",x"C0",x"06", -- 0x0338
    x"03",x"60",x"06",x"03",x"80",x"02",x"04",x"A0", -- 0x0340
    x"04",x"03",x"E0",x"02",x"02",x"A0",x"02",x"05", -- 0x0348
    x"E0",x"02",x"04",x"C0",x"02",x"04",x"60",x"08", -- 0x0350
    x"02",x"A0",x"04",x"03",x"80",x"0C",x"01",x"E0", -- 0x0358
    x"06",x"02",x"80",x"06",x"03",x"80",x"02",x"04", -- 0x0360
    x"80",x"04",x"04",x"C0",x"02",x"03",x"E0",x"02", -- 0x0368
    x"04",x"A0",x"02",x"04",x"E0",x"02",x"04",x"60", -- 0x0370
    x"08",x"01",x"E0",x"04",x"03",x"80",x"0C",x"01", -- 0x0378
    x"A0",x"06",x"02",x"E0",x"06",x"02",x"80",x"02", -- 0x0380
    x"04",x"60",x"04",x"03",x"A0",x"02",x"04",x"80", -- 0x0388
    x"02",x"05",x"C0",x"02",x"04",x"A0",x"02",x"05", -- 0x0390
    x"3A",x"D6",x"83",x"3D",x"C0",x"3A",x"9B",x"82", -- 0x0398
    x"A7",x"C0",x"32",x"B4",x"83",x"CD",x"DD",x"0A", -- 0x03A0
    x"CD",x"3C",x"06",x"CD",x"C6",x"32",x"AF",x"32", -- 0x03A8
    x"5B",x"82",x"CD",x"DB",x"29",x"21",x"50",x"A8", -- 0x03B0
    x"CD",x"6B",x"2A",x"CD",x"CD",x"09",x"CD",x"23", -- 0x03B8
    x"20",x"3E",x"01",x"32",x"5B",x"82",x"32",x"9B", -- 0x03C0
    x"82",x"C9",x"3A",x"D6",x"83",x"3D",x"C0",x"3A", -- 0x03C8
    x"9B",x"82",x"A7",x"C8",x"CD",x"F6",x"33",x"CD", -- 0x03D0
    x"DE",x"2A",x"CD",x"40",x"34",x"CD",x"65",x"09", -- 0x03D8
    x"CD",x"93",x"08",x"CD",x"8E",x"30",x"CD",x"8B", -- 0x03E0
    x"28",x"CD",x"48",x"22",x"CD",x"81",x"27",x"CD", -- 0x03E8
    x"50",x"30",x"CD",x"40",x"25",x"C9",x"3A",x"6C", -- 0x03F0
    x"82",x"B7",x"C0",x"3A",x"04",x"80",x"A7",x"C0", -- 0x03F8
    x"3A",x"99",x"82",x"A7",x"C2",x"6F",x"34",x"11", -- 0x0400
    x"47",x"80",x"3E",x"30",x"32",x"99",x"82",x"21", -- 0x0408
    x"9A",x"82",x"34",x"4E",x"06",x"00",x"21",x"3E", -- 0x0410
    x"0F",x"09",x"4E",x"0C",x"CA",x"35",x"34",x"21", -- 0x0418
    x"25",x"34",x"09",x"E5",x"21",x"44",x"80",x"C9", -- 0x0420
    x"C3",x"29",x"2D",x"C3",x"CA",x"2C",x"C3",x"6D", -- 0x0428
    x"2C",x"C3",x"14",x"2C",x"C9",x"AF",x"32",x"9A", -- 0x0430
    x"82",x"32",x"99",x"82",x"32",x"5B",x"82",x"C9", -- 0x0438
    x"21",x"44",x"80",x"11",x"47",x"80",x"3A",x"48", -- 0x0440
    x"82",x"A7",x"C2",x"43",x"2C",x"32",x"4C",x"82", -- 0x0448
    x"3A",x"49",x"82",x"A7",x"C2",x"96",x"2C",x"32", -- 0x0450
    x"4D",x"82",x"3A",x"4A",x"82",x"A7",x"C2",x"FF", -- 0x0458
    x"2C",x"32",x"4E",x"82",x"3A",x"4B",x"82",x"A7", -- 0x0460
    x"C2",x"5E",x"2D",x"32",x"4F",x"82",x"C9",x"3D", -- 0x0468
    x"32",x"99",x"82",x"C9",x"3A",x"23",x"81",x"3C", -- 0x0470
    x"32",x"23",x"81",x"FE",x"06",x"D8",x"AF",x"32", -- 0x0478
    x"23",x"81",x"C9",x"3A",x"FD",x"83",x"4F",x"3A", -- 0x0480
    x"23",x"81",x"32",x"21",x"81",x"FE",x"01",x"CA", -- 0x0488
    x"A7",x"34",x"FE",x"02",x"CA",x"BC",x"34",x"FE", -- 0x0490
    x"03",x"CA",x"D1",x"34",x"FE",x"04",x"CA",x"E6", -- 0x0498
    x"34",x"FE",x"05",x"CA",x"FB",x"34",x"C9",x"0D", -- 0x04A0
    x"20",x"0B",x"3A",x"5E",x"82",x"A7",x"C0",x"21", -- 0x04A8
    x"64",x"AB",x"C3",x"10",x"35",x"3A",x"63",x"82", -- 0x04B0
    x"A7",x"C0",x"18",x"F3",x"0D",x"20",x"0B",x"3A", -- 0x04B8
    x"5F",x"82",x"A7",x"C0",x"21",x"A4",x"AA",x"C3", -- 0x04C0
    x"10",x"35",x"3A",x"64",x"82",x"A7",x"C0",x"18", -- 0x04C8
    x"F3",x"0D",x"20",x"0B",x"3A",x"60",x"82",x"A7", -- 0x04D0
    x"C0",x"21",x"E4",x"A9",x"C3",x"10",x"35",x"3A", -- 0x04D8
    x"65",x"82",x"A7",x"C0",x"18",x"F3",x"0D",x"20", -- 0x04E0
    x"0B",x"3A",x"61",x"82",x"A7",x"C0",x"21",x"24", -- 0x04E8
    x"A9",x"C3",x"10",x"35",x"3A",x"66",x"82",x"A7", -- 0x04F0
    x"C0",x"18",x"F3",x"0D",x"20",x"0B",x"3A",x"62", -- 0x04F8
    x"82",x"A7",x"C0",x"21",x"64",x"A8",x"C3",x"10", -- 0x0500
    x"35",x"3A",x"67",x"82",x"A7",x"C0",x"18",x"F3", -- 0x0508
    x"36",x"2C",x"23",x"36",x"2D",x"01",x"1F",x"00", -- 0x0510
    x"09",x"36",x"2E",x"23",x"36",x"2F",x"C9",x"3A", -- 0x0518
    x"FD",x"83",x"4F",x"3A",x"23",x"81",x"32",x"20", -- 0x0520
    x"81",x"FE",x"01",x"CA",x"43",x"35",x"FE",x"02", -- 0x0528
    x"CA",x"58",x"35",x"FE",x"03",x"CA",x"6D",x"35", -- 0x0530
    x"FE",x"04",x"CA",x"82",x"35",x"FE",x"05",x"CA", -- 0x0538
    x"97",x"35",x"C9",x"0D",x"20",x"0B",x"3A",x"5E", -- 0x0540
    x"82",x"A7",x"C0",x"21",x"64",x"AB",x"C3",x"AC", -- 0x0548
    x"35",x"3A",x"63",x"82",x"A7",x"C0",x"18",x"F3", -- 0x0550
    x"0D",x"20",x"0B",x"3A",x"5F",x"82",x"A7",x"C0", -- 0x0558
    x"21",x"A4",x"AA",x"C3",x"AC",x"35",x"3A",x"64", -- 0x0560
    x"82",x"A7",x"C0",x"18",x"F3",x"0D",x"20",x"0B", -- 0x0568
    x"3A",x"60",x"82",x"A7",x"C0",x"21",x"E4",x"A9", -- 0x0570
    x"C3",x"AC",x"35",x"3A",x"65",x"82",x"A7",x"C0", -- 0x0578
    x"18",x"F3",x"0D",x"20",x"0B",x"3A",x"61",x"82", -- 0x0580
    x"A7",x"C0",x"21",x"24",x"A9",x"C3",x"AC",x"35", -- 0x0588
    x"3A",x"66",x"82",x"A7",x"C0",x"18",x"F3",x"0D", -- 0x0590
    x"20",x"0B",x"3A",x"62",x"82",x"A7",x"C0",x"21", -- 0x0598
    x"64",x"A8",x"C3",x"AC",x"35",x"3A",x"67",x"82", -- 0x05A0
    x"A7",x"C0",x"18",x"F3",x"36",x"10",x"23",x"36", -- 0x05A8
    x"10",x"01",x"1F",x"00",x"09",x"36",x"D0",x"23", -- 0x05B0
    x"36",x"D1",x"C9",x"3A",x"FD",x"83",x"4F",x"3A", -- 0x05B8
    x"20",x"81",x"32",x"21",x"81",x"FE",x"01",x"CA", -- 0x05C0
    x"DF",x"35",x"FE",x"02",x"CA",x"F4",x"35",x"FE", -- 0x05C8
    x"03",x"CA",x"09",x"36",x"FE",x"04",x"CA",x"1E", -- 0x05D0
    x"36",x"FE",x"05",x"CA",x"33",x"36",x"C9",x"0D", -- 0x05D8
    x"20",x"0B",x"3A",x"5E",x"82",x"A7",x"C0",x"21", -- 0x05E0
    x"64",x"AB",x"C3",x"48",x"36",x"3A",x"63",x"82", -- 0x05E8
    x"A7",x"C0",x"18",x"F3",x"0D",x"20",x"0B",x"3A", -- 0x05F0
    x"5F",x"82",x"A7",x"C0",x"21",x"A4",x"AA",x"C3", -- 0x05F8
    x"48",x"36",x"3A",x"64",x"82",x"A7",x"C0",x"18", -- 0x0600
    x"F3",x"0D",x"20",x"0B",x"3A",x"60",x"82",x"A7", -- 0x0608
    x"C0",x"21",x"E4",x"A9",x"C3",x"48",x"36",x"3A", -- 0x0610
    x"65",x"82",x"A7",x"C0",x"18",x"F3",x"0D",x"20", -- 0x0618
    x"0B",x"3A",x"61",x"82",x"A7",x"C0",x"21",x"24", -- 0x0620
    x"A9",x"C3",x"48",x"36",x"3A",x"66",x"82",x"A7", -- 0x0628
    x"C0",x"18",x"F3",x"0D",x"20",x"0B",x"3A",x"62", -- 0x0630
    x"82",x"A7",x"C0",x"21",x"64",x"A8",x"C3",x"48", -- 0x0638
    x"36",x"3A",x"67",x"82",x"A7",x"C0",x"18",x"F3", -- 0x0640
    x"36",x"D0",x"23",x"36",x"D1",x"01",x"1F",x"00", -- 0x0648
    x"09",x"36",x"D2",x"23",x"36",x"D3",x"C9",x"3A", -- 0x0650
    x"FD",x"83",x"4F",x"3A",x"21",x"81",x"FE",x"01", -- 0x0658
    x"CA",x"78",x"36",x"FE",x"02",x"CA",x"8D",x"36", -- 0x0660
    x"FE",x"03",x"CA",x"A2",x"36",x"FE",x"04",x"CA", -- 0x0668
    x"B7",x"36",x"FE",x"05",x"CA",x"CC",x"36",x"C9", -- 0x0670
    x"0D",x"20",x"0B",x"3A",x"5E",x"82",x"A7",x"C0", -- 0x0678
    x"21",x"64",x"AB",x"C3",x"E1",x"36",x"3A",x"63", -- 0x0680
    x"82",x"A7",x"C0",x"18",x"F3",x"0D",x"20",x"0B", -- 0x0688
    x"3A",x"5F",x"82",x"A7",x"C0",x"21",x"A4",x"AA", -- 0x0690
    x"C3",x"E1",x"36",x"3A",x"64",x"82",x"A7",x"C0", -- 0x0698
    x"18",x"F3",x"0D",x"20",x"0B",x"3A",x"60",x"82", -- 0x06A0
    x"A7",x"C0",x"21",x"E4",x"A9",x"C3",x"E1",x"36", -- 0x06A8
    x"3A",x"65",x"82",x"A7",x"C0",x"18",x"F3",x"0D", -- 0x06B0
    x"20",x"0B",x"3A",x"61",x"82",x"A7",x"C0",x"21", -- 0x06B8
    x"24",x"A9",x"C3",x"E1",x"36",x"3A",x"66",x"82", -- 0x06C0
    x"A7",x"C0",x"18",x"F3",x"0D",x"20",x"0B",x"3A", -- 0x06C8
    x"62",x"82",x"A7",x"C0",x"21",x"64",x"A8",x"C3", -- 0x06D0
    x"E1",x"36",x"3A",x"67",x"82",x"A7",x"C0",x"18", -- 0x06D8
    x"F3",x"36",x"10",x"23",x"36",x"10",x"01",x"1F", -- 0x06E0
    x"00",x"09",x"36",x"10",x"23",x"36",x"10",x"3A", -- 0x06E8
    x"04",x"80",x"A7",x"C0",x"AF",x"32",x"21",x"81", -- 0x06F0
    x"32",x"20",x"81",x"C9",x"3A",x"20",x"81",x"A7", -- 0x06F8
    x"C2",x"1C",x"37",x"21",x"5C",x"80",x"70",x"23", -- 0x0700
    x"36",x"19",x"23",x"36",x"03",x"23",x"36",x"20", -- 0x0708
    x"3E",x"A0",x"32",x"40",x"83",x"11",x"20",x"00", -- 0x0710
    x"CD",x"03",x"09",x"C9",x"3E",x"01",x"32",x"04", -- 0x0718
    x"80",x"E1",x"C9",x"21",x"5C",x"80",x"AF",x"77", -- 0x0720
    x"23",x"77",x"23",x"77",x"23",x"77",x"C9",x"3A", -- 0x0728
    x"34",x"81",x"A7",x"C2",x"79",x"37",x"DD",x"21", -- 0x0730
    x"1B",x"81",x"DD",x"7E",x"01",x"A7",x"CC",x"96", -- 0x0738
    x"37",x"3A",x"3D",x"81",x"CB",x"47",x"C2",x"3C", -- 0x0740
    x"38",x"3A",x"35",x"81",x"A7",x"20",x"01",x"C9", -- 0x0748
    x"3A",x"34",x"81",x"A7",x"20",x"23",x"CD",x"B8", -- 0x0750
    x"37",x"3A",x"47",x"80",x"FE",x"5A",x"D8",x"FE", -- 0x0758
    x"68",x"D0",x"3A",x"40",x"80",x"47",x"3A",x"44", -- 0x0760
    x"80",x"C6",x"04",x"B8",x"D8",x"D6",x"08",x"B8", -- 0x0768
    x"D0",x"3E",x"01",x"32",x"34",x"81",x"3E",x"18", -- 0x0770
    x"DF",x"DD",x"21",x"44",x"80",x"FD",x"21",x"40", -- 0x0778
    x"80",x"DD",x"7E",x"00",x"FD",x"77",x"00",x"DD", -- 0x0780
    x"7E",x"01",x"FD",x"77",x"01",x"DD",x"7E",x"03", -- 0x0788
    x"C6",x"02",x"FD",x"77",x"03",x"C9",x"3A",x"35", -- 0x0790
    x"81",x"A7",x"C0",x"21",x"3D",x"81",x"34",x"21", -- 0x0798
    x"41",x"80",x"36",x"1E",x"23",x"36",x"04",x"23", -- 0x07A0
    x"36",x"60",x"3E",x"01",x"32",x"35",x"81",x"32", -- 0x07A8
    x"3D",x"83",x"3E",x"3C",x"32",x"3E",x"83",x"C9", -- 0x07B0
    x"21",x"3E",x"83",x"7E",x"A7",x"28",x"2B",x"35", -- 0x07B8
    x"3E",x"3C",x"CB",x"3F",x"BE",x"20",x"0F",x"2B", -- 0x07C0
    x"7E",x"A7",x"3E",x"21",x"32",x"41",x"80",x"F0", -- 0x07C8
    x"3E",x"A1",x"32",x"41",x"80",x"C9",x"2B",x"7E", -- 0x07D0
    x"E6",x"7F",x"21",x"28",x"38",x"3C",x"CD",x"23", -- 0x07D8
    x"38",x"7E",x"21",x"1C",x"81",x"86",x"32",x"40", -- 0x07E0
    x"80",x"C9",x"2B",x"7E",x"A7",x"F2",x"F2",x"37", -- 0x07E8
    x"35",x"35",x"34",x"7E",x"E6",x"7F",x"21",x"28", -- 0x07F0
    x"38",x"CD",x"23",x"38",x"7E",x"FE",x"01",x"38", -- 0x07F8
    x"0A",x"28",x"1A",x"21",x"1C",x"81",x"86",x"32", -- 0x0800
    x"40",x"80",x"C9",x"21",x"3D",x"83",x"7E",x"EE", -- 0x0808
    x"80",x"77",x"3E",x"3C",x"32",x"3E",x"83",x"3E", -- 0x0810
    x"1E",x"32",x"41",x"80",x"C9",x"3E",x"3C",x"32", -- 0x0818
    x"3E",x"83",x"C9",x"85",x"6F",x"D0",x"24",x"C9", -- 0x0820
    x"00",x"EE",x"EC",x"EA",x"E8",x"E6",x"E4",x"E2", -- 0x0828
    x"E0",x"01",x"DE",x"DC",x"DA",x"D8",x"D6",x"D4", -- 0x0830
    x"D2",x"D0",x"00",x"D0",x"3A",x"35",x"81",x"A7", -- 0x0838
    x"C8",x"AF",x"32",x"34",x"81",x"21",x"40",x"80", -- 0x0840
    x"AF",x"77",x"23",x"77",x"23",x"77",x"23",x"77", -- 0x0848
    x"32",x"35",x"81",x"C9",x"21",x"40",x"80",x"70", -- 0x0850
    x"23",x"36",x"19",x"23",x"36",x"03",x"23",x"36", -- 0x0858
    x"10",x"3E",x"A0",x"32",x"40",x"83",x"C9",x"21", -- 0x0860
    x"40",x"80",x"AF",x"77",x"23",x"77",x"23",x"77", -- 0x0868
    x"23",x"77",x"C9",x"3A",x"B7",x"83",x"FE",x"02", -- 0x0870
    x"DA",x"FC",x"38",x"FE",x"05",x"D2",x"FD",x"38", -- 0x0878
    x"3A",x"01",x"81",x"A7",x"CC",x"15",x"39",x"3A", -- 0x0880
    x"4F",x"81",x"A7",x"C8",x"21",x"46",x"81",x"7E", -- 0x0888
    x"23",x"BE",x"C2",x"39",x"39",x"35",x"11",x"06", -- 0x0890
    x"A8",x"3A",x"50",x"81",x"CB",x"47",x"CA",x"F6", -- 0x0898
    x"38",x"21",x"9C",x"24",x"AF",x"47",x"3A",x"4E", -- 0x08A0
    x"81",x"4F",x"3C",x"3C",x"32",x"4E",x"81",x"09", -- 0x08A8
    x"06",x"00",x"EB",x"3A",x"45",x"81",x"4F",x"09", -- 0x08B0
    x"EB",x"0E",x"20",x"3A",x"45",x"81",x"81",x"32", -- 0x08B8
    x"45",x"81",x"7E",x"12",x"23",x"13",x"7E",x"12", -- 0x08C0
    x"3A",x"4E",x"81",x"FE",x"10",x"D8",x"AF",x"32", -- 0x08C8
    x"4F",x"81",x"32",x"4E",x"81",x"32",x"45",x"81", -- 0x08D0
    x"32",x"46",x"81",x"32",x"47",x"81",x"C9",x"3A", -- 0x08D8
    x"FE",x"83",x"FE",x"02",x"C0",x"AF",x"32",x"4F", -- 0x08E0
    x"81",x"32",x"4E",x"81",x"32",x"45",x"81",x"32", -- 0x08E8
    x"46",x"81",x"32",x"47",x"81",x"C9",x"21",x"8C", -- 0x08F0
    x"24",x"C3",x"A4",x"38",x"C9",x"3A",x"01",x"81", -- 0x08F8
    x"A7",x"CC",x"07",x"39",x"C3",x"87",x"38",x"3A", -- 0x0900
    x"4F",x"81",x"A7",x"C0",x"3E",x"01",x"32",x"50", -- 0x0908
    x"81",x"CD",x"25",x"39",x"C9",x"3A",x"4F",x"81", -- 0x0910
    x"A7",x"C0",x"3A",x"50",x"81",x"3C",x"32",x"50", -- 0x0918
    x"81",x"CD",x"25",x"39",x"C9",x"3A",x"9B",x"81", -- 0x0920
    x"E6",x"0F",x"87",x"87",x"87",x"21",x"46",x"81", -- 0x0928
    x"77",x"23",x"77",x"3E",x"01",x"32",x"4F",x"81", -- 0x0930
    x"C9",x"7E",x"A7",x"28",x"02",x"35",x"C9",x"3A", -- 0x0938
    x"46",x"81",x"77",x"C9",x"3A",x"50",x"81",x"CB", -- 0x0940
    x"47",x"C8",x"3A",x"B7",x"83",x"FE",x"02",x"D8", -- 0x0948
    x"3A",x"47",x"80",x"C6",x"08",x"FE",x"2A",x"D8", -- 0x0950
    x"FE",x"3B",x"D0",x"3A",x"44",x"80",x"C6",x"08", -- 0x0958
    x"47",x"3A",x"01",x"81",x"4F",x"C6",x"08",x"B8", -- 0x0960
    x"D8",x"79",x"D6",x"20",x"B8",x"D0",x"79",x"D6", -- 0x0968
    x"08",x"B8",x"30",x"04",x"CD",x"59",x"23",x"C9", -- 0x0970
    x"3E",x"01",x"32",x"04",x"80",x"21",x"46",x"A8", -- 0x0978
    x"36",x"68",x"23",x"36",x"69",x"01",x"1F",x"00", -- 0x0980
    x"09",x"36",x"6A",x"23",x"36",x"6B",x"C9",x"3A", -- 0x0988
    x"FE",x"83",x"A7",x"C8",x"3A",x"A2",x"81",x"FE", -- 0x0990
    x"0F",x"D0",x"FE",x"02",x"D8",x"3A",x"40",x"81", -- 0x0998
    x"A7",x"C0",x"3E",x"D0",x"DF",x"C9",x"3A",x"01", -- 0x09A0
    x"81",x"A7",x"20",x"05",x"AF",x"32",x"3F",x"83", -- 0x09A8
    x"C9",x"3A",x"50",x"81",x"CB",x"47",x"C8",x"3A", -- 0x09B0
    x"4F",x"81",x"A7",x"C0",x"21",x"3F",x"83",x"34", -- 0x09B8
    x"7E",x"FE",x"40",x"28",x"05",x"FE",x"70",x"28", -- 0x09C0
    x"13",x"C9",x"21",x"46",x"A8",x"36",x"68",x"23", -- 0x09C8
    x"36",x"69",x"01",x"1F",x"00",x"09",x"36",x"6A", -- 0x09D0
    x"23",x"36",x"6B",x"C9",x"21",x"46",x"A8",x"36", -- 0x09D8
    x"D0",x"23",x"36",x"D1",x"01",x"1F",x"00",x"09", -- 0x09E0
    x"36",x"D2",x"23",x"36",x"D3",x"AF",x"32",x"3F", -- 0x09E8
    x"83",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DF8
    x"21",x"E2",x"83",x"7E",x"B7",x"3A",x"00",x"E0", -- 0x0E00
    x"2F",x"20",x"04",x"E6",x"C4",x"77",x"C9",x"E6", -- 0x0E08
    x"C4",x"C0",x"3C",x"CD",x"A7",x"07",x"AF",x"32", -- 0x0E10
    x"86",x"83",x"ED",x"5B",x"D4",x"83",x"CB",x"76", -- 0x0E18
    x"C2",x"3E",x"3E",x"CB",x"56",x"77",x"20",x"09", -- 0x0E20
    x"3C",x"32",x"18",x"B8",x"3E",x"04",x"32",x"7E", -- 0x0E28
    x"83",x"21",x"36",x"3E",x"19",x"E9",x"18",x"24", -- 0x0E30
    x"18",x"1B",x"18",x"19",x"18",x"1E",x"77",x"3C", -- 0x0E38
    x"32",x"1C",x"B8",x"3E",x"04",x"32",x"7F",x"83", -- 0x0E40
    x"21",x"4D",x"3E",x"19",x"E9",x"18",x"0D",x"18", -- 0x0E48
    x"04",x"18",x"11",x"18",x"13",x"21",x"E3",x"83", -- 0x0E50
    x"34",x"CB",x"46",x"C0",x"0E",x"01",x"18",x"0A", -- 0x0E58
    x"0E",x"02",x"18",x"06",x"0E",x"03",x"18",x"02", -- 0x0E60
    x"0E",x"06",x"3A",x"E1",x"83",x"81",x"27",x"30", -- 0x0E68
    x"02",x"3E",x"99",x"32",x"E1",x"83",x"3A",x"FE", -- 0x0E70
    x"83",x"B7",x"C0",x"3A",x"D6",x"83",x"FE",x"05", -- 0x0E78
    x"CC",x"13",x"0D",x"3E",x"05",x"32",x"D6",x"83", -- 0x0E80
    x"AF",x"32",x"D8",x"83",x"21",x"40",x"80",x"11", -- 0x0E88
    x"41",x"80",x"01",x"1F",x"00",x"70",x"ED",x"B0", -- 0x0E90
    x"C3",x"8A",x"0B",x"21",x"D8",x"83",x"36",x"FF", -- 0x0E98
    x"CD",x"79",x"07",x"AF",x"32",x"9B",x"82",x"32", -- 0x0EA0
    x"21",x"80",x"3E",x"05",x"32",x"1B",x"80",x"3E", -- 0x0EA8
    x"03",x"32",x"2B",x"80",x"11",x"F2",x"0F",x"21", -- 0x0EB0
    x"8D",x"AA",x"06",x"0B",x"EF",x"3A",x"E4",x"83", -- 0x0EB8
    x"FE",x"0A",x"D0",x"21",x"15",x"AB",x"CD",x"CC", -- 0x0EC0
    x"0B",x"11",x"3F",x"10",x"06",x"07",x"EF",x"11", -- 0x0EC8
    x"09",x"10",x"06",x"04",x"EF",x"11",x"28",x"10", -- 0x0ED0
    x"06",x"07",x"EF",x"C9",x"FF",x"FF",x"FF",x"FF", -- 0x0ED8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F00
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F08
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F10
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F18
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F20
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F28
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F40
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F48
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F50
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F58
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F60
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F68
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F70
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
