-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_PGM_23 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_PGM_23 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"0B",x"06",x"FF",x"1E",x"0C",x"FF",x"C9",x"21", -- 0x0000
    x"40",x"45",x"35",x"C0",x"2C",x"34",x"21",x"3D", -- 0x0008
    x"0F",x"CD",x"AD",x"0E",x"11",x"86",x"06",x"FF", -- 0x0010
    x"11",x"92",x"06",x"FF",x"11",x"8B",x"06",x"FF", -- 0x0018
    x"11",x"8C",x"06",x"FF",x"11",x"00",x"02",x"FF", -- 0x0020
    x"C9",x"21",x"40",x"45",x"35",x"C0",x"21",x"02", -- 0x0028
    x"48",x"22",x"0B",x"40",x"21",x"09",x"40",x"36", -- 0x0030
    x"20",x"21",x"41",x"45",x"34",x"C9",x"2A",x"0B", -- 0x0038
    x"40",x"06",x"1A",x"3E",x"10",x"D7",x"11",x"06", -- 0x0040
    x"00",x"19",x"22",x"0B",x"40",x"21",x"09",x"40", -- 0x0048
    x"35",x"C0",x"21",x"1D",x"0F",x"CD",x"AD",x"0E", -- 0x0050
    x"11",x"0D",x"06",x"FF",x"21",x"81",x"10",x"11", -- 0x0058
    x"60",x"40",x"01",x"18",x"00",x"ED",x"B0",x"21", -- 0x0060
    x"99",x"10",x"22",x"44",x"45",x"21",x"4A",x"4A", -- 0x0068
    x"22",x"46",x"45",x"21",x"40",x"45",x"36",x"32", -- 0x0070
    x"2C",x"34",x"2C",x"36",x"0B",x"2C",x"36",x"06", -- 0x0078
    x"C9",x"50",x"1C",x"00",x"4A",x"50",x"1E",x"00", -- 0x0080
    x"62",x"50",x"1A",x"06",x"7B",x"50",x"10",x"04", -- 0x0088
    x"92",x"50",x"26",x"05",x"A9",x"50",x"33",x"01", -- 0x0090
    x"C2",x"0C",x"0C",x"0C",x"10",x"10",x"05",x"00", -- 0x0098
    x"10",x"20",x"24",x"23",x"0C",x"0C",x"0C",x"10", -- 0x00A0
    x"10",x"08",x"00",x"10",x"20",x"24",x"23",x"0C", -- 0x00A8
    x"0C",x"0C",x"10",x"01",x"00",x"00",x"10",x"20", -- 0x00B0
    x"24",x"23",x"0C",x"0C",x"0C",x"10",x"01",x"05", -- 0x00B8
    x"00",x"10",x"20",x"24",x"23",x"0C",x"0C",x"0C", -- 0x00C0
    x"10",x"08",x"00",x"00",x"10",x"20",x"24",x"23", -- 0x00C8
    x"0C",x"0C",x"0C",x"10",x"1D",x"29",x"23",x"24", -- 0x00D0
    x"15",x"22",x"29",x"21",x"40",x"45",x"35",x"C0", -- 0x00D8
    x"36",x"05",x"2A",x"44",x"45",x"7E",x"23",x"22", -- 0x00E0
    x"44",x"45",x"2A",x"46",x"45",x"77",x"11",x"E0", -- 0x00E8
    x"FF",x"19",x"22",x"46",x"45",x"21",x"42",x"45", -- 0x00F0
    x"35",x"C0",x"36",x"0B",x"21",x"40",x"45",x"36", -- 0x00F8
    x"14",x"2C",x"34",x"C9",x"21",x"40",x"45",x"35", -- 0x0100
    x"C0",x"36",x"01",x"2C",x"35",x"2A",x"46",x"45", -- 0x0108
    x"11",x"63",x"01",x"19",x"22",x"46",x"45",x"21", -- 0x0110
    x"43",x"45",x"35",x"C0",x"21",x"40",x"45",x"36", -- 0x0118
    x"96",x"2C",x"34",x"34",x"C9",x"21",x"40",x"45", -- 0x0120
    x"35",x"C0",x"2C",x"34",x"21",x"60",x"40",x"3E", -- 0x0128
    x"10",x"06",x"18",x"D7",x"CD",x"F6",x"18",x"CD", -- 0x0130
    x"17",x"19",x"21",x"BD",x"0E",x"C3",x"AD",x"0E", -- 0x0138
    x"21",x"41",x"45",x"34",x"CD",x"CF",x"12",x"CD", -- 0x0140
    x"F5",x"13",x"3E",x"01",x"32",x"19",x"40",x"21", -- 0x0148
    x"01",x"00",x"22",x"80",x"43",x"22",x"A0",x"43", -- 0x0150
    x"AF",x"32",x"82",x"43",x"32",x"0D",x"40",x"21", -- 0x0158
    x"00",x"41",x"06",x"40",x"D7",x"21",x"B5",x"31", -- 0x0160
    x"11",x"18",x"41",x"7E",x"12",x"23",x"13",x"7E", -- 0x0168
    x"12",x"23",x"7E",x"32",x"1D",x"41",x"11",x"02", -- 0x0170
    x"07",x"FF",x"3E",x"20",x"32",x"15",x"41",x"21", -- 0x0178
    x"05",x"41",x"36",x"FF",x"2C",x"36",x"05",x"11", -- 0x0180
    x"07",x"06",x"FF",x"C9",x"CD",x"4B",x"1B",x"CD", -- 0x0188
    x"37",x"25",x"CD",x"38",x"26",x"CD",x"AA",x"2A", -- 0x0190
    x"CD",x"C0",x"2F",x"21",x"80",x"43",x"7E",x"2C", -- 0x0198
    x"B6",x"0F",x"D8",x"21",x"41",x"45",x"36",x"00", -- 0x01A0
    x"C9",x"3A",x"02",x"40",x"A7",x"C8",x"21",x"05", -- 0x01A8
    x"40",x"34",x"AF",x"32",x"0A",x"40",x"C9",x"21", -- 0x01B0
    x"47",x"12",x"E5",x"3A",x"0A",x"40",x"EF",x"C5", -- 0x01B8
    x"11",x"F3",x"11",x"39",x"12",x"AF",x"32",x"19", -- 0x01C0
    x"40",x"3E",x"01",x"32",x"04",x"68",x"3D",x"32", -- 0x01C8
    x"03",x"68",x"21",x"DD",x"0E",x"CD",x"AD",x"0E", -- 0x01D0
    x"21",x"60",x"40",x"06",x"40",x"AF",x"D7",x"32", -- 0x01D8
    x"B0",x"40",x"32",x"06",x"40",x"21",x"02",x"48", -- 0x01E0
    x"22",x"0B",x"40",x"21",x"09",x"40",x"36",x"10", -- 0x01E8
    x"2C",x"34",x"C9",x"2A",x"0B",x"40",x"06",x"1D", -- 0x01F0
    x"3E",x"10",x"D7",x"11",x"03",x"00",x"19",x"06", -- 0x01F8
    x"1D",x"D7",x"19",x"22",x"0B",x"40",x"21",x"09", -- 0x0200
    x"40",x"35",x"C0",x"2C",x"34",x"AF",x"32",x"06", -- 0x0208
    x"68",x"32",x"07",x"68",x"32",x"0D",x"40",x"11", -- 0x0210
    x"01",x"07",x"FF",x"11",x"01",x"06",x"FF",x"1E", -- 0x0218
    x"16",x"FF",x"1C",x"FF",x"3A",x"17",x"40",x"47", -- 0x0220
    x"E6",x"0F",x"32",x"78",x"49",x"78",x"E6",x"F0", -- 0x0228
    x"C8",x"0F",x"0F",x"0F",x"0F",x"32",x"98",x"49", -- 0x0230
    x"C9",x"3A",x"02",x"40",x"A7",x"C8",x"3D",x"11", -- 0x0238
    x"18",x"06",x"28",x"01",x"1C",x"FF",x"C9",x"3A", -- 0x0240
    x"11",x"40",x"CB",x"7F",x"C2",x"87",x"12",x"CB", -- 0x0248
    x"77",x"C8",x"3A",x"02",x"40",x"FE",x"02",x"D8", -- 0x0250
    x"D6",x"02",x"32",x"02",x"40",x"21",x"00",x"01", -- 0x0258
    x"22",x"0D",x"40",x"AF",x"32",x"0A",x"40",x"3E", -- 0x0260
    x"03",x"32",x"05",x"40",x"3E",x"01",x"32",x"06", -- 0x0268
    x"40",x"11",x"04",x"06",x"FF",x"CD",x"9D",x"12", -- 0x0270
    x"CD",x"0E",x"31",x"11",x"00",x"04",x"FF",x"3A", -- 0x0278
    x"0E",x"40",x"0F",x"D0",x"1C",x"FF",x"C9",x"3A", -- 0x0280
    x"02",x"40",x"A7",x"28",x"0A",x"3D",x"32",x"02", -- 0x0288
    x"40",x"21",x"00",x"00",x"C3",x"60",x"12",x"3E", -- 0x0290
    x"01",x"32",x"05",x"40",x"C9",x"AF",x"21",x"00", -- 0x0298
    x"41",x"47",x"D7",x"21",x"30",x"42",x"06",x"10", -- 0x02A0
    x"D7",x"21",x"60",x"40",x"06",x"40",x"D7",x"21", -- 0x02A8
    x"60",x"42",x"01",x"02",x"B0",x"DF",x"32",x"19", -- 0x02B0
    x"40",x"21",x"00",x"41",x"11",x"01",x"41",x"01", -- 0x02B8
    x"C0",x"00",x"36",x"00",x"ED",x"B0",x"3A",x"07", -- 0x02C0
    x"40",x"32",x"48",x"41",x"32",x"88",x"41",x"21", -- 0x02C8
    x"C0",x"41",x"11",x"28",x"C9",x"06",x"20",x"72", -- 0x02D0
    x"2C",x"73",x"2C",x"10",x"FA",x"C9",x"3A",x"0A", -- 0x02D8
    x"40",x"EF",x"0E",x"13",x"30",x"13",x"48",x"13", -- 0x02E0
    x"D2",x"13",x"FF",x"17",x"62",x"18",x"B1",x"18", -- 0x02E8
    x"3F",x"19",x"03",x"1A",x"7A",x"1A",x"3A",x"0A", -- 0x02F0
    x"40",x"EF",x"0E",x"13",x"30",x"13",x"8D",x"13", -- 0x02F8
    x"D2",x"13",x"FF",x"17",x"62",x"18",x"8E",x"19", -- 0x0300
    x"C4",x"19",x"03",x"1A",x"7A",x"1A",x"AF",x"32", -- 0x0308
    x"19",x"40",x"21",x"60",x"40",x"06",x"40",x"D7", -- 0x0310
    x"21",x"0A",x"40",x"34",x"2D",x"36",x"20",x"21", -- 0x0318
    x"00",x"48",x"22",x"0B",x"40",x"CD",x"17",x"19", -- 0x0320
    x"3E",x"01",x"32",x"06",x"40",x"C3",x"CF",x"12", -- 0x0328
    x"2A",x"0B",x"40",x"06",x"20",x"3E",x"10",x"D7", -- 0x0330
    x"22",x"0B",x"40",x"21",x"09",x"40",x"35",x"C0", -- 0x0338
    x"2C",x"34",x"21",x"BD",x"0E",x"C3",x"AD",x"0E", -- 0x0340
    x"AF",x"32",x"5F",x"42",x"32",x"06",x"68",x"32", -- 0x0348
    x"07",x"68",x"32",x"0D",x"40",x"21",x"0A",x"40", -- 0x0350
    x"34",x"2D",x"36",x"96",x"3A",x"0E",x"40",x"0F", -- 0x0358
    x"38",x"25",x"11",x"00",x"05",x"FF",x"1E",x"02", -- 0x0360
    x"FF",x"14",x"FF",x"1E",x"04",x"FF",x"11",x"03", -- 0x0368
    x"07",x"FF",x"1E",x"00",x"FF",x"21",x"40",x"41", -- 0x0370
    x"11",x"00",x"41",x"01",x"40",x"00",x"ED",x"B0", -- 0x0378
    x"2A",x"1D",x"41",x"22",x"18",x"41",x"C9",x"11", -- 0x0380
    x"01",x"05",x"FF",x"18",x"D5",x"AF",x"32",x"5F", -- 0x0388
    x"42",x"3A",x"0F",x"40",x"0F",x"30",x"08",x"3E", -- 0x0390
    x"01",x"32",x"06",x"68",x"32",x"07",x"68",x"3E", -- 0x0398
    x"01",x"32",x"0D",x"40",x"21",x"0A",x"40",x"34", -- 0x03A0
    x"2D",x"36",x"96",x"11",x"00",x"05",x"FF",x"1C", -- 0x03A8
    x"FF",x"1C",x"FF",x"11",x"03",x"06",x"FF",x"1C", -- 0x03B0
    x"FF",x"11",x"03",x"07",x"FF",x"1E",x"00",x"FF", -- 0x03B8
    x"21",x"80",x"41",x"11",x"00",x"41",x"01",x"40", -- 0x03C0
    x"00",x"ED",x"B0",x"2A",x"1D",x"41",x"22",x"18", -- 0x03C8
    x"41",x"C9",x"21",x"09",x"40",x"35",x"C0",x"36", -- 0x03D0
    x"20",x"2C",x"34",x"11",x"82",x"06",x"FF",x"1E", -- 0x03D8
    x"07",x"FF",x"CD",x"F6",x"18",x"CD",x"17",x"19", -- 0x03E0
    x"CD",x"CF",x"12",x"AF",x"32",x"19",x"40",x"21", -- 0x03E8
    x"60",x"40",x"06",x"40",x"D7",x"21",x"19",x"48", -- 0x03F0
    x"11",x"1C",x"00",x"06",x"1E",x"3E",x"36",x"0E", -- 0x03F8
    x"39",x"77",x"2C",x"71",x"2C",x"71",x"2C",x"71", -- 0x0400
    x"2C",x"71",x"19",x"10",x"F4",x"C9",x"C8",x"2E", -- 0x0408
    x"D0",x"36",x"28",x"63",x"28",x"5E",x"00",x"D0", -- 0x0410
    x"36",x"D0",x"2D",x"28",x"5E",x"30",x"63",x"00", -- 0x0418
    x"D8",x"36",x"D8",x"36",x"30",x"5E",x"30",x"5E", -- 0x0420
    x"02",x"D8",x"2F",x"E0",x"36",x"38",x"63",x"38", -- 0x0428
    x"5E",x"00",x"E0",x"36",x"D8",x"31",x"38",x"5E", -- 0x0430
    x"40",x"63",x"00",x"D0",x"30",x"C8",x"30",x"48", -- 0x0438
    x"62",x"48",x"62",x"00",x"C0",x"30",x"B8",x"31", -- 0x0440
    x"48",x"5D",x"50",x"62",x"00",x"B8",x"36",x"B8", -- 0x0448
    x"35",x"50",x"5E",x"5F",x"62",x"00",x"B0",x"34", -- 0x0450
    x"B8",x"2C",x"5F",x"5D",x"5F",x"60",x"00",x"C0", -- 0x0458
    x"35",x"B8",x"34",x"50",x"60",x"48",x"60",x"00", -- 0x0460
    x"C0",x"2D",x"C8",x"2C",x"48",x"62",x"50",x"62", -- 0x0468
    x"00",x"D0",x"36",x"D0",x"2C",x"50",x"60",x"50", -- 0x0470
    x"62",x"00",x"D8",x"2D",x"D8",x"31",x"5F",x"62", -- 0x0478
    x"5F",x"60",x"00",x"D0",x"32",x"C8",x"31",x"5F", -- 0x0480
    x"62",x"5F",x"60",x"00",x"C0",x"32",x"C0",x"2F", -- 0x0488
    x"50",x"60",x"48",x"60",x"00",x"C8",x"2F",x"C8", -- 0x0490
    x"33",x"48",x"62",x"48",x"60",x"00",x"C8",x"2C", -- 0x0498
    x"D0",x"2C",x"40",x"60",x"38",x"60",x"00",x"D0", -- 0x04A0
    x"30",x"D0",x"2D",x"38",x"62",x"40",x"62",x"00", -- 0x04A8
    x"D0",x"31",x"C8",x"34",x"48",x"62",x"48",x"60", -- 0x04B0
    x"00",x"C8",x"30",x"C0",x"30",x"40",x"60",x"38", -- 0x04B8
    x"61",x"00",x"B8",x"30",x"B0",x"30",x"38",x"62", -- 0x04C0
    x"40",x"63",x"00",x"B0",x"2C",x"B0",x"30",x"40", -- 0x04C8
    x"60",x"38",x"61",x"00",x"B0",x"36",x"B0",x"2C", -- 0x04D0
    x"30",x"60",x"30",x"62",x"00",x"B8",x"2C",x"B8", -- 0x04D8
    x"30",x"38",x"62",x"38",x"60",x"00",x"B8",x"2C", -- 0x04E0
    x"C0",x"2C",x"30",x"60",x"30",x"62",x"00",x"C8", -- 0x04E8
    x"36",x"C0",x"30",x"38",x"62",x"40",x"5C",x"00", -- 0x04F0
    x"C0",x"2C",x"C8",x"35",x"38",x"60",x"30",x"61", -- 0x04F8
    x"00",x"C0",x"30",x"C0",x"2C",x"28",x"5E",x"28", -- 0x0500
    x"60",x"00",x"C0",x"31",x"B8",x"30",x"28",x"62", -- 0x0508
    x"30",x"62",x"00",x"B0",x"32",x"B0",x"36",x"38", -- 0x0510
    x"62",x"40",x"62",x"00",x"B0",x"2E",x"B8",x"2D", -- 0x0518
    x"48",x"62",x"50",x"62",x"00",x"C0",x"2E",x"C8", -- 0x0520
    x"2D",x"5F",x"62",x"5F",x"3A",x"00",x"D0",x"36", -- 0x0528
    x"D0",x"36",x"5F",x"3A",x"5F",x"60",x"01",x"D0", -- 0x0530
    x"36",x"D0",x"36",x"50",x"3A",x"50",x"3A",x"02", -- 0x0538
    x"D0",x"36",x"D0",x"36",x"5F",x"62",x"5F",x"3A", -- 0x0540
    x"01",x"D0",x"36",x"D0",x"36",x"5F",x"3A",x"5F", -- 0x0548
    x"3A",x"02",x"D0",x"36",x"D0",x"2E",x"5F",x"3A", -- 0x0550
    x"5F",x"3A",x"00",x"D8",x"36",x"D8",x"36",x"5F", -- 0x0558
    x"3A",x"5F",x"60",x"04",x"D8",x"36",x"D8",x"36", -- 0x0560
    x"50",x"60",x"48",x"60",x"04",x"D0",x"32",x"D0", -- 0x0568
    x"36",x"40",x"60",x"38",x"60",x"00",x"D0",x"36", -- 0x0570
    x"D0",x"36",x"30",x"3A",x"30",x"3A",x"01",x"C8", -- 0x0578
    x"31",x"C0",x"32",x"30",x"3A",x"30",x"3A",x"00", -- 0x0580
    x"C0",x"36",x"C0",x"36",x"30",x"3A",x"30",x"3A", -- 0x0588
    x"01",x"B8",x"31",x"B0",x"32",x"30",x"3A",x"30", -- 0x0590
    x"60",x"00",x"B0",x"36",x"B0",x"36",x"28",x"3A", -- 0x0598
    x"28",x"3A",x"00",x"B0",x"36",x"B0",x"36",x"28", -- 0x05A0
    x"3A",x"28",x"3A",x"00",x"B0",x"2E",x"B8",x"2D", -- 0x05A8
    x"30",x"62",x"30",x"3A",x"00",x"C0",x"36",x"C0", -- 0x05B0
    x"2E",x"30",x"3A",x"30",x"3A",x"00",x"C8",x"36", -- 0x05B8
    x"C8",x"36",x"38",x"62",x"40",x"62",x"04",x"C8", -- 0x05C0
    x"36",x"C8",x"36",x"48",x"62",x"48",x"3A",x"01", -- 0x05C8
    x"C8",x"2E",x"D0",x"36",x"48",x"3A",x"50",x"62", -- 0x05D0
    x"00",x"D0",x"36",x"D0",x"36",x"5F",x"62",x"5F", -- 0x05D8
    x"3A",x"04",x"D0",x"36",x"D0",x"2D",x"5F",x"3A", -- 0x05E0
    x"5F",x"60",x"00",x"D8",x"36",x"D8",x"36",x"50", -- 0x05E8
    x"60",x"48",x"60",x"01",x"D8",x"36",x"D8",x"36", -- 0x05F0
    x"40",x"60",x"38",x"60",x"02",x"D0",x"31",x"C8", -- 0x05F8
    x"32",x"30",x"60",x"28",x"60",x"00",x"C0",x"31", -- 0x0600
    x"B8",x"30",x"28",x"62",x"30",x"62",x"00",x"B0", -- 0x0608
    x"32",x"B0",x"36",x"38",x"62",x"40",x"62",x"00", -- 0x0610
    x"B0",x"2E",x"B8",x"2D",x"48",x"62",x"50",x"62", -- 0x0618
    x"00",x"C0",x"2E",x"C8",x"2D",x"5F",x"62",x"5F", -- 0x0620
    x"3A",x"00",x"D0",x"36",x"D0",x"36",x"5F",x"3A", -- 0x0628
    x"5F",x"60",x"01",x"D0",x"36",x"D0",x"36",x"50", -- 0x0630
    x"3A",x"50",x"3A",x"01",x"D0",x"36",x"D0",x"36", -- 0x0638
    x"5F",x"62",x"5F",x"3A",x"02",x"D0",x"36",x"D0", -- 0x0640
    x"36",x"5F",x"3A",x"5F",x"3A",x"02",x"D0",x"36", -- 0x0648
    x"D0",x"2E",x"5F",x"3A",x"5F",x"3A",x"00",x"D8", -- 0x0650
    x"36",x"D8",x"36",x"5F",x"3A",x"5F",x"60",x"01", -- 0x0658
    x"D8",x"36",x"D8",x"36",x"50",x"60",x"48",x"60", -- 0x0660
    x"01",x"D0",x"32",x"D0",x"36",x"40",x"60",x"38", -- 0x0668
    x"60",x"00",x"D0",x"36",x"D0",x"36",x"30",x"3A", -- 0x0670
    x"30",x"3A",x"04",x"C8",x"31",x"C0",x"32",x"30", -- 0x0678
    x"3A",x"30",x"3A",x"00",x"C0",x"36",x"C0",x"36", -- 0x0680
    x"30",x"3A",x"30",x"3A",x"01",x"B8",x"31",x"B0", -- 0x0688
    x"32",x"30",x"3A",x"30",x"60",x"00",x"B0",x"36", -- 0x0690
    x"B0",x"36",x"28",x"3A",x"28",x"3A",x"00",x"B0", -- 0x0698
    x"36",x"B0",x"36",x"28",x"3A",x"28",x"3A",x"00", -- 0x06A0
    x"B0",x"2E",x"B8",x"2D",x"30",x"62",x"30",x"3A", -- 0x06A8
    x"00",x"C0",x"36",x"C0",x"2E",x"30",x"3A",x"30", -- 0x06B0
    x"3A",x"00",x"C8",x"36",x"C8",x"36",x"38",x"62", -- 0x06B8
    x"40",x"62",x"04",x"C8",x"36",x"C8",x"36",x"48", -- 0x06C0
    x"62",x"48",x"3A",x"04",x"C8",x"2E",x"D0",x"36", -- 0x06C8
    x"48",x"3A",x"50",x"62",x"00",x"D0",x"36",x"D0", -- 0x06D0
    x"36",x"5F",x"62",x"5F",x"3A",x"01",x"D0",x"36", -- 0x06D8
    x"D0",x"2D",x"5F",x"3A",x"5F",x"60",x"00",x"D8", -- 0x06E0
    x"36",x"D8",x"36",x"50",x"60",x"48",x"60",x"04", -- 0x06E8
    x"D8",x"36",x"D8",x"36",x"40",x"60",x"38",x"60", -- 0x06F0
    x"04",x"D0",x"31",x"C8",x"32",x"30",x"60",x"28", -- 0x06F8
    x"60",x"00",x"C8",x"2C",x"D0",x"2C",x"28",x"62", -- 0x0700
    x"30",x"62",x"00",x"D8",x"2C",x"E0",x"36",x"38", -- 0x0708
    x"62",x"40",x"62",x"00",x"E0",x"36",x"E0",x"36", -- 0x0710
    x"48",x"62",x"50",x"62",x"01",x"E0",x"36",x"D8", -- 0x0718
    x"34",x"5F",x"5C",x"50",x"60",x"00",x"E0",x"36", -- 0x0720
    x"E0",x"36",x"48",x"60",x"40",x"60",x"02",x"E0", -- 0x0728
    x"36",x"E0",x"36",x"38",x"60",x"30",x"60",x"01", -- 0x0730
    x"E0",x"36",x"E0",x"36",x"28",x"5E",x"30",x"62", -- 0x0738
    x"01",x"D8",x"34",x"E0",x"36",x"36",x"5C",x"30", -- 0x0740
    x"60",x"00",x"E0",x"36",x"E0",x"36",x"28",x"5E", -- 0x0748
    x"30",x"5C",x"04",x"E0",x"36",x"E0",x"36",x"28", -- 0x0750
    x"5E",x"30",x"62",x"01",x"E0",x"36",x"E0",x"36", -- 0x0758
    x"38",x"62",x"40",x"62",x"04",x"D8",x"30",x"D0", -- 0x0760
    x"30",x"48",x"62",x"57",x"5C",x"00",x"C8",x"30", -- 0x0768
    x"C0",x"30",x"48",x"60",x"40",x"60",x"00",x"B8", -- 0x0770
    x"30",x"B0",x"34",x"38",x"60",x"30",x"60",x"00", -- 0x0778
    x"B8",x"2C",x"C0",x"2C",x"28",x"3A",x"28",x"3A", -- 0x0780
    x"00",x"C8",x"2C",x"D0",x"2C",x"28",x"3A",x"28", -- 0x0788
    x"3A",x"00",x"D8",x"2C",x"D8",x"34",x"28",x"3A", -- 0x0790
    x"28",x"3A",x"00",x"E0",x"36",x"E0",x"36",x"28", -- 0x0798
    x"3A",x"30",x"5C",x"01",x"E0",x"36",x"E0",x"36", -- 0x07A0
    x"28",x"3A",x"28",x"3A",x"02",x"D8",x"30",x"D0", -- 0x07A8
    x"34",x"28",x"3A",x"28",x"3A",x"00",x"D8",x"2C", -- 0x07B0
    x"E0",x"36",x"28",x"3A",x"28",x"3A",x"00",x"E0", -- 0x07B8
    x"36",x"E0",x"36",x"28",x"3A",x"28",x"3A",x"01", -- 0x07C0
    x"E0",x"36",x"E0",x"36",x"28",x"3A",x"28",x"3A", -- 0x07C8
    x"01",x"E0",x"36",x"E0",x"36",x"28",x"3A",x"28", -- 0x07D0
    x"3A",x"01",x"E0",x"36",x"D8",x"34",x"28",x"3A", -- 0x07D8
    x"28",x"3A",x"00",x"E0",x"36",x"E0",x"36",x"28", -- 0x07E0
    x"3A",x"28",x"3A",x"04",x"E0",x"36",x"D8",x"30", -- 0x07E8
    x"28",x"3A",x"28",x"3A",x"00",x"D0",x"30",x"C8", -- 0x07F0
    x"30",x"28",x"3A",x"28",x"60",x"00",x"FF",x"21", -- 0x07F8
    x"09",x"40",x"35",x"C0",x"36",x"0A",x"2C",x"34", -- 0x0800
    x"3E",x"01",x"32",x"19",x"40",x"21",x"01",x"00", -- 0x0808
    x"22",x"80",x"43",x"22",x"A0",x"43",x"AF",x"32", -- 0x0810
    x"82",x"43",x"21",x"08",x"41",x"35",x"11",x"03", -- 0x0818
    x"07",x"FF",x"21",x"10",x"41",x"11",x"11",x"41", -- 0x0820
    x"01",x"0D",x"00",x"36",x"00",x"ED",x"B0",x"21", -- 0x0828
    x"B5",x"31",x"3A",x"1E",x"41",x"47",x"87",x"80", -- 0x0830
    x"5F",x"16",x"00",x"19",x"7E",x"32",x"18",x"41", -- 0x0838
    x"23",x"7E",x"32",x"19",x"41",x"23",x"7E",x"32", -- 0x0840
    x"1D",x"41",x"11",x"02",x"07",x"FF",x"3E",x"08", -- 0x0848
    x"32",x"15",x"41",x"3E",x"FF",x"32",x"05",x"41", -- 0x0850
    x"3E",x"05",x"32",x"06",x"41",x"11",x"00",x"07", -- 0x0858
    x"FF",x"C9",x"CD",x"4B",x"1B",x"CD",x"37",x"25", -- 0x0860
    x"CD",x"38",x"26",x"CD",x"AA",x"2A",x"CD",x"C0", -- 0x0868
    x"2F",x"CD",x"1B",x"1B",x"CD",x"7B",x"31",x"CD", -- 0x0870
    x"26",x"1B",x"21",x"80",x"43",x"7E",x"0F",x"38", -- 0x0878
    x"19",x"2C",x"7E",x"0F",x"D8",x"21",x"80",x"43", -- 0x0880
    x"11",x"81",x"43",x"36",x"00",x"01",x"A0",x"01", -- 0x0888
    x"ED",x"B0",x"21",x"0A",x"40",x"34",x"2D",x"36", -- 0x0890
    x"64",x"C9",x"3A",x"12",x"41",x"FE",x"FF",x"C0", -- 0x0898
    x"21",x"80",x"45",x"36",x"96",x"2C",x"36",x"00", -- 0x08A0
    x"21",x"0A",x"40",x"36",x"08",x"2D",x"36",x"64", -- 0x08A8
    x"C9",x"3A",x"08",x"41",x"A7",x"20",x"28",x"CD", -- 0x08B0
    x"F6",x"18",x"CD",x"17",x"19",x"11",x"00",x"06", -- 0x08B8
    x"FF",x"1E",x"02",x"FF",x"3E",x"01",x"32",x"04", -- 0x08C0
    x"68",x"3D",x"32",x"03",x"68",x"21",x"C0",x"45", -- 0x08C8
    x"36",x"96",x"2C",x"36",x"00",x"3E",x"09",x"32", -- 0x08D0
    x"0A",x"40",x"AF",x"32",x"19",x"40",x"C9",x"3A", -- 0x08D8
    x"0E",x"40",x"0F",x"38",x"09",x"21",x"0A",x"40", -- 0x08E0
    x"36",x"03",x"2D",x"36",x"32",x"C9",x"21",x"0A", -- 0x08E8
    x"40",x"34",x"2D",x"36",x"32",x"C9",x"21",x"03", -- 0x08F0
    x"48",x"11",x"05",x"00",x"0E",x"20",x"3E",x"10", -- 0x08F8
    x"06",x"1B",x"77",x"23",x"10",x"FC",x"19",x"0D", -- 0x0900
    x"20",x"F6",x"21",x"2A",x"40",x"06",x"19",x"AF", -- 0x0908
    x"77",x"2C",x"77",x"2C",x"10",x"FA",x"C9",x"21", -- 0x0910
    x"80",x"42",x"11",x"81",x"42",x"01",x"A0",x"02", -- 0x0918
    x"36",x"00",x"ED",x"B0",x"21",x"60",x"42",x"11", -- 0x0920
    x"61",x"42",x"01",x"1F",x"00",x"36",x"00",x"ED", -- 0x0928
    x"B0",x"21",x"60",x"40",x"11",x"61",x"40",x"01", -- 0x0930
    x"3F",x"00",x"36",x"00",x"ED",x"B0",x"C9",x"21", -- 0x0938
    x"09",x"40",x"35",x"C0",x"3A",x"08",x"41",x"A7", -- 0x0940
    x"20",x"10",x"3A",x"0E",x"40",x"0F",x"38",x"19", -- 0x0948
    x"3E",x"01",x"32",x"05",x"40",x"AF",x"32",x"41", -- 0x0950
    x"45",x"C9",x"3A",x"88",x"41",x"A7",x"20",x"19", -- 0x0958
    x"21",x"0A",x"40",x"36",x"03",x"2D",x"36",x"01", -- 0x0960
    x"C9",x"3A",x"88",x"41",x"A7",x"20",x"0A",x"3E", -- 0x0968
    x"01",x"32",x"05",x"40",x"AF",x"32",x"41",x"45", -- 0x0970
    x"C9",x"21",x"00",x"41",x"11",x"40",x"41",x"01", -- 0x0978
    x"40",x"00",x"ED",x"B0",x"AF",x"32",x"0A",x"40", -- 0x0980
    x"3E",x"04",x"32",x"05",x"40",x"C9",x"3A",x"08", -- 0x0988
    x"41",x"A7",x"20",x"28",x"CD",x"F6",x"18",x"CD", -- 0x0990
    x"17",x"19",x"11",x"00",x"06",x"FF",x"1E",x"03", -- 0x0998
    x"FF",x"3E",x"01",x"32",x"04",x"68",x"3D",x"32", -- 0x09A0
    x"03",x"68",x"21",x"C0",x"45",x"36",x"96",x"2C", -- 0x09A8
    x"36",x"00",x"3E",x"09",x"32",x"0A",x"40",x"AF", -- 0x09B0
    x"32",x"19",x"40",x"C9",x"21",x"0A",x"40",x"34", -- 0x09B8
    x"2D",x"36",x"64",x"C9",x"21",x"09",x"40",x"35", -- 0x09C0
    x"C0",x"3A",x"08",x"41",x"A7",x"20",x"10",x"3A", -- 0x09C8
    x"48",x"41",x"A7",x"20",x"0A",x"3E",x"01",x"32", -- 0x09D0
    x"05",x"40",x"AF",x"32",x"41",x"45",x"C9",x"3A", -- 0x09D8
    x"48",x"41",x"A7",x"20",x"09",x"21",x"0A",x"40", -- 0x09E0
    x"36",x"03",x"2D",x"36",x"01",x"C9",x"21",x"00", -- 0x09E8
    x"41",x"11",x"80",x"41",x"01",x"40",x"00",x"ED", -- 0x09F0
    x"B0",x"AF",x"32",x"0A",x"40",x"3E",x"03",x"32", -- 0x09F8
    x"05",x"40",x"C9",x"3A",x"81",x"45",x"EF",x"0D", -- 0x0A00
    x"1A",x"35",x"1A",x"50",x"1A",x"CD",x"4B",x"1B", -- 0x0A08
    x"CD",x"37",x"25",x"CD",x"38",x"26",x"CD",x"C0", -- 0x0A10
    x"2F",x"21",x"80",x"45",x"35",x"C0",x"36",x"05", -- 0x0A18
    x"2C",x"34",x"3E",x"01",x"32",x"04",x"68",x"3E", -- 0x0A20
    x"00",x"32",x"03",x"68",x"32",x"19",x"40",x"3E", -- 0x0A28
    x"08",x"32",x"02",x"82",x"C9",x"21",x"80",x"45", -- 0x0A30
    x"35",x"C0",x"2C",x"34",x"CD",x"F6",x"18",x"11", -- 0x0A38
    x"08",x"06",x"FF",x"1C",x"FF",x"1C",x"FF",x"21", -- 0x0A40
    x"5D",x"0F",x"CD",x"AD",x"0E",x"C3",x"17",x"19", -- 0x0A48
    x"21",x"80",x"45",x"35",x"C0",x"21",x"08",x"41", -- 0x0A50
    x"34",x"21",x"00",x"41",x"34",x"11",x"00",x"07", -- 0x0A58
    x"FF",x"AF",x"32",x"5F",x"42",x"21",x"0A",x"40", -- 0x0A60
    x"36",x"03",x"2D",x"36",x"0A",x"CD",x"CF",x"12", -- 0x0A68
    x"AF",x"32",x"1E",x"41",x"21",x"BD",x"0E",x"C3", -- 0x0A70
    x"AD",x"0E",x"3A",x"C1",x"45",x"EF",x"84",x"1A", -- 0x0A78
    x"98",x"1A",x"B7",x"1A",x"21",x"C0",x"45",x"35", -- 0x0A80
    x"C0",x"2C",x"34",x"11",x"80",x"06",x"FF",x"1E", -- 0x0A88
    x"82",x"FF",x"21",x"3D",x"0F",x"C3",x"AD",x"0E", -- 0x0A90
    x"CD",x"C5",x"1A",x"7D",x"FE",x"0A",x"28",x"0B", -- 0x0A98
    x"87",x"87",x"5F",x"16",x"00",x"21",x"2F",x"40", -- 0x0AA0
    x"19",x"36",x"00",x"11",x"00",x"02",x"FF",x"21", -- 0x0AA8
    x"C0",x"45",x"36",x"80",x"2C",x"34",x"C9",x"21", -- 0x0AB0
    x"C0",x"45",x"35",x"C0",x"21",x"0A",x"40",x"36", -- 0x0AB8
    x"07",x"2D",x"36",x"64",x"C9",x"01",x"1E",x"00", -- 0x0AC0
    x"11",x"03",x"00",x"6A",x"DD",x"21",x"A2",x"40", -- 0x0AC8
    x"3A",x"0D",x"40",x"0F",x"30",x"02",x"DD",x"19", -- 0x0AD0
    x"FD",x"21",x"00",x"42",x"DD",x"7E",x"02",x"FD", -- 0x0AD8
    x"BE",x"02",x"20",x"0F",x"DD",x"7E",x"01",x"FD", -- 0x0AE0
    x"BE",x"01",x"20",x"07",x"DD",x"7E",x"00",x"FD", -- 0x0AE8
    x"BE",x"00",x"C8",x"30",x"09",x"FD",x"19",x"2C", -- 0x0AF0
    x"0D",x"0D",x"0D",x"C8",x"18",x"DE",x"7D",x"21", -- 0x0AF8
    x"1D",x"42",x"11",x"20",x"42",x"ED",x"B8",x"6F", -- 0x0B00
    x"DD",x"7E",x"00",x"FD",x"77",x"00",x"DD",x"7E", -- 0x0B08
    x"01",x"FD",x"77",x"01",x"DD",x"7E",x"02",x"FD", -- 0x0B10
    x"77",x"02",x"C9",x"3A",x"5F",x"42",x"E6",x"3F", -- 0x0B18
    x"C0",x"11",x"0C",x"03",x"FF",x"C9",x"3A",x"07", -- 0x0B20
    x"41",x"A7",x"C0",x"21",x"A4",x"40",x"3A",x"0D", -- 0x0B28
    x"40",x"0F",x"30",x"03",x"21",x"A7",x"40",x"7E", -- 0x0B30
    x"A7",x"C8",x"CD",x"B0",x"31",x"21",x"08",x"41", -- 0x0B38
    x"34",x"11",x"03",x"07",x"FF",x"3E",x"01",x"32", -- 0x0B40
    x"07",x"41",x"C9",x"CD",x"24",x"1D",x"CD",x"36", -- 0x0B48
    x"20",x"CD",x"4F",x"1E",x"CD",x"97",x"21",x"CD", -- 0x0B50
    x"BF",x"22",x"CD",x"89",x"23",x"CD",x"C8",x"24", -- 0x0B58
    x"C3",x"29",x"1E",x"DD",x"7E",x"0E",x"A7",x"28", -- 0x0B60
    x"05",x"3D",x"DD",x"77",x"0E",x"C9",x"DD",x"6E", -- 0x0B68
    x"0C",x"DD",x"66",x"0D",x"7E",x"FE",x"FF",x"28", -- 0x0B70
    x"15",x"DD",x"77",x"16",x"23",x"7E",x"DD",x"77", -- 0x0B78
    x"12",x"23",x"7E",x"DD",x"77",x"0E",x"23",x"DD", -- 0x0B80
    x"75",x"0C",x"DD",x"74",x"0D",x"C9",x"23",x"7E", -- 0x0B88
    x"DD",x"77",x"0C",x"23",x"7E",x"DD",x"77",x"0D", -- 0x0B90
    x"18",x"C9",x"DD",x"E5",x"E1",x"3E",x"07",x"85", -- 0x0B98
    x"6F",x"DD",x"36",x"0A",x"00",x"DD",x"7E",x"05", -- 0x0BA0
    x"DD",x"BE",x"03",x"28",x"04",x"38",x"1E",x"18", -- 0x0BA8
    x"56",x"DD",x"7E",x"06",x"DD",x"BE",x"04",x"28", -- 0x0BB0
    x"0E",x"38",x"06",x"36",x"00",x"2C",x"36",x"01", -- 0x0BB8
    x"C9",x"36",x"00",x"2C",x"36",x"FF",x"C9",x"36", -- 0x0BC0
    x"00",x"2C",x"36",x"00",x"C9",x"DD",x"7E",x"06", -- 0x0BC8
    x"DD",x"BE",x"04",x"28",x"2C",x"38",x"15",x"36", -- 0x0BD0
    x"FF",x"2C",x"36",x"01",x"DD",x"7E",x"03",x"DD", -- 0x0BD8
    x"96",x"05",x"47",x"DD",x"7E",x"06",x"DD",x"96", -- 0x0BE0
    x"04",x"4F",x"18",x"55",x"36",x"FF",x"2C",x"36", -- 0x0BE8
    x"FF",x"DD",x"7E",x"03",x"DD",x"96",x"05",x"47", -- 0x0BF0
    x"DD",x"7E",x"04",x"DD",x"96",x"06",x"4F",x"18", -- 0x0BF8
    x"40",x"36",x"FF",x"2C",x"36",x"00",x"C9",x"DD", -- 0x0C00
    x"7E",x"06",x"DD",x"BE",x"04",x"28",x"2C",x"38", -- 0x0C08
    x"15",x"36",x"01",x"2C",x"36",x"01",x"DD",x"7E", -- 0x0C10
    x"05",x"DD",x"96",x"03",x"47",x"DD",x"7E",x"06", -- 0x0C18
    x"DD",x"96",x"04",x"4F",x"18",x"1B",x"36",x"01", -- 0x0C20
    x"2C",x"36",x"FF",x"DD",x"7E",x"05",x"DD",x"96", -- 0x0C28
    x"03",x"47",x"DD",x"7E",x"04",x"DD",x"96",x"06", -- 0x0C30
    x"4F",x"18",x"06",x"36",x"01",x"2C",x"36",x"00", -- 0x0C38
    x"C9",x"79",x"B8",x"28",x"16",x"38",x"0B",x"DD", -- 0x0C40
    x"36",x"09",x"00",x"CD",x"64",x"1C",x"DD",x"77", -- 0x0C48
    x"0B",x"C9",x"DD",x"36",x"09",x"01",x"78",x"41", -- 0x0C50
    x"4F",x"18",x"F0",x"DD",x"36",x"09",x"01",x"DD", -- 0x0C58
    x"36",x"0B",x"FF",x"C9",x"AF",x"67",x"68",x"57", -- 0x0C60
    x"59",x"06",x"08",x"CB",x"FF",x"07",x"29",x"A7", -- 0x0C68
    x"ED",x"52",x"38",x"03",x"10",x"F5",x"C9",x"19", -- 0x0C70
    x"CB",x"87",x"10",x"EF",x"C9",x"DD",x"7E",x"04", -- 0x0C78
    x"DD",x"BE",x"06",x"28",x"4A",x"DD",x"7E",x"03", -- 0x0C80
    x"DD",x"BE",x"05",x"28",x"58",x"DD",x"CB",x"09", -- 0x0C88
    x"46",x"28",x"1E",x"DD",x"7E",x"07",x"DD",x"86", -- 0x0C90
    x"03",x"DD",x"77",x"03",x"DD",x"7E",x"0B",x"DD", -- 0x0C98
    x"86",x"0A",x"DD",x"77",x"0A",x"D0",x"DD",x"7E", -- 0x0CA0
    x"08",x"DD",x"86",x"04",x"DD",x"77",x"04",x"A7", -- 0x0CA8
    x"C9",x"DD",x"7E",x"08",x"DD",x"86",x"04",x"DD", -- 0x0CB0
    x"77",x"04",x"DD",x"7E",x"0B",x"DD",x"86",x"0A", -- 0x0CB8
    x"DD",x"77",x"0A",x"D0",x"DD",x"7E",x"07",x"DD", -- 0x0CC0
    x"86",x"03",x"DD",x"77",x"03",x"A7",x"C9",x"DD", -- 0x0CC8
    x"7E",x"03",x"DD",x"BE",x"05",x"28",x"0C",x"30", -- 0x0CD0
    x"05",x"DD",x"34",x"03",x"A7",x"C9",x"DD",x"35", -- 0x0CD8
    x"03",x"A7",x"C9",x"37",x"C9",x"DD",x"7E",x"04", -- 0x0CE0
    x"DD",x"BE",x"06",x"30",x"05",x"DD",x"34",x"04", -- 0x0CE8
    x"A7",x"C9",x"DD",x"35",x"04",x"A7",x"C9",x"DD", -- 0x0CF0
    x"6E",x"13",x"DD",x"66",x"14",x"7E",x"FE",x"80", -- 0x0CF8
    x"20",x"0C",x"23",x"7E",x"DD",x"77",x"13",x"23", -- 0x0D00
    x"7E",x"DD",x"77",x"14",x"18",x"E9",x"DD",x"86", -- 0x0D08
    x"03",x"DD",x"77",x"03",x"23",x"7E",x"DD",x"86", -- 0x0D10
    x"04",x"DD",x"77",x"04",x"23",x"DD",x"75",x"13", -- 0x0D18
    x"DD",x"74",x"14",x"C9",x"DD",x"21",x"10",x"41", -- 0x0D20
    x"DD",x"7E",x"05",x"A7",x"20",x"12",x"DD",x"7E", -- 0x0D28
    x"04",x"DD",x"77",x"05",x"DD",x"7E",x"06",x"E6", -- 0x0D30
    x"0F",x"CC",x"44",x"1D",x"DD",x"34",x"06",x"C9", -- 0x0D38
    x"DD",x"35",x"05",x"C9",x"CD",x"4A",x"1D",x"C3", -- 0x0D40
    x"D8",x"1D",x"FD",x"2A",x"18",x"41",x"3E",x"01", -- 0x0D48
    x"32",x"10",x"41",x"32",x"30",x"42",x"DD",x"7E", -- 0x0D50
    x"06",x"2F",x"E6",x"F0",x"47",x"6F",x"26",x"12", -- 0x0D58
    x"29",x"29",x"E5",x"FD",x"7E",x"02",x"E6",x"F8", -- 0x0D60
    x"0F",x"0F",x"0F",x"5F",x"16",x"00",x"19",x"22", -- 0x0D68
    x"35",x"42",x"FD",x"7E",x"03",x"32",x"34",x"42", -- 0x0D70
    x"E1",x"1E",x"20",x"19",x"FD",x"7E",x"00",x"E6", -- 0x0D78
    x"F8",x"0F",x"0F",x"0F",x"5F",x"19",x"22",x"32", -- 0x0D80
    x"42",x"FD",x"7E",x"01",x"32",x"31",x"42",x"78", -- 0x0D88
    x"0F",x"0F",x"5F",x"21",x"C0",x"41",x"19",x"FD", -- 0x0D90
    x"7E",x"02",x"77",x"2C",x"36",x"28",x"2C",x"FD", -- 0x0D98
    x"7E",x"00",x"77",x"2C",x"36",x"28",x"AF",x"32", -- 0x0DA0
    x"38",x"42",x"32",x"11",x"41",x"2A",x"18",x"41", -- 0x0DA8
    x"1E",x"09",x"FD",x"7E",x"04",x"A7",x"20",x"02", -- 0x0DB0
    x"1E",x"06",x"19",x"22",x"18",x"41",x"FD",x"7E", -- 0x0DB8
    x"04",x"A7",x"28",x"05",x"FD",x"7E",x"08",x"18", -- 0x0DC0
    x"03",x"FD",x"7E",x"05",x"32",x"1A",x"41",x"2A", -- 0x0DC8
    x"35",x"42",x"2B",x"2B",x"22",x"1B",x"41",x"C9", -- 0x0DD0
    x"FD",x"7E",x"04",x"A7",x"C8",x"68",x"26",x"12", -- 0x0DD8
    x"29",x"29",x"E5",x"FD",x"7E",x"06",x"E6",x"F8", -- 0x0DE0
    x"0F",x"0F",x"0F",x"5F",x"19",x"22",x"3D",x"42", -- 0x0DE8
    x"FD",x"7E",x"07",x"32",x"3C",x"42",x"E1",x"1E", -- 0x0DF0
    x"20",x"19",x"FD",x"7E",x"04",x"E6",x"F8",x"0F", -- 0x0DF8
    x"0F",x"0F",x"5F",x"19",x"22",x"3A",x"42",x"FD", -- 0x0E00
    x"7E",x"05",x"32",x"39",x"42",x"78",x"0F",x"0F", -- 0x0E08
    x"5F",x"21",x"C0",x"41",x"19",x"2C",x"FD",x"7E", -- 0x0E10
    x"06",x"77",x"2C",x"2C",x"FD",x"7E",x"04",x"77", -- 0x0E18
    x"3E",x"01",x"32",x"11",x"41",x"32",x"38",x"42", -- 0x0E20
    x"C9",x"DD",x"21",x"00",x"45",x"11",x"03",x"00", -- 0x0E28
    x"06",x"04",x"CD",x"3A",x"1E",x"DD",x"19",x"10", -- 0x0E30
    x"F9",x"C9",x"DD",x"CB",x"00",x"46",x"C8",x"DD", -- 0x0E38
    x"7E",x"02",x"D6",x"03",x"DD",x"77",x"02",x"FE", -- 0x0E40
    x"1F",x"D0",x"DD",x"CB",x"00",x"86",x"C9",x"DD", -- 0x0E48
    x"21",x"80",x"43",x"DD",x"7E",x"00",x"DD",x"B6", -- 0x0E50
    x"01",x"0F",x"D0",x"DD",x"7E",x"02",x"EF",x"73", -- 0x0E58
    x"1E",x"9A",x"1E",x"5C",x"1F",x"8F",x"1F",x"90", -- 0x0E60
    x"1F",x"91",x"1F",x"92",x"1F",x"AD",x"1F",x"E6", -- 0x0E68
    x"1F",x"E7",x"1F",x"DD",x"36",x"03",x"58",x"DD", -- 0x0E70
    x"36",x"23",x"58",x"DD",x"36",x"04",x"D0",x"DD", -- 0x0E78
    x"36",x"24",x"E0",x"21",x"E8",x"1F",x"22",x"8C", -- 0x0E80
    x"43",x"21",x"F7",x"1F",x"22",x"AC",x"43",x"DD", -- 0x0E88
    x"36",x"0E",x"00",x"DD",x"36",x"2E",x"00",x"DD", -- 0x0E90
    x"34",x"02",x"21",x"06",x"41",x"35",x"20",x"1B", -- 0x0E98
    x"3A",x"00",x"41",x"A7",x"28",x"07",x"3D",x"28", -- 0x0EA0
    x"08",x"36",x"04",x"18",x"06",x"36",x"06",x"18", -- 0x0EA8
    x"02",x"36",x"05",x"2D",x"35",x"20",x"04",x"DD", -- 0x0EB0
    x"34",x"02",x"C9",x"DD",x"21",x"A0",x"43",x"CD", -- 0x0EB8
    x"63",x"1B",x"DD",x"21",x"80",x"43",x"CD",x"63", -- 0x0EC0
    x"1B",x"CD",x"CF",x"1E",x"C3",x"25",x"1F",x"3A", -- 0x0EC8
    x"06",x"40",x"0F",x"30",x"1B",x"3A",x"0D",x"40", -- 0x0ED0
    x"0F",x"38",x"33",x"3A",x"12",x"40",x"06",x"00", -- 0x0ED8
    x"CB",x"67",x"28",x"02",x"CB",x"C0",x"CB",x"77", -- 0x0EE0
    x"28",x"02",x"CB",x"C8",x"78",x"0F",x"30",x"0E", -- 0x0EE8
    x"DD",x"7E",x"03",x"3D",x"FE",x"38",x"D8",x"DD", -- 0x0EF0
    x"77",x"03",x"DD",x"35",x"23",x"C9",x"0F",x"D0", -- 0x0EF8
    x"DD",x"7E",x"03",x"3C",x"FE",x"D8",x"D0",x"DD", -- 0x0F00
    x"77",x"03",x"DD",x"34",x"23",x"C9",x"3A",x"12", -- 0x0F08
    x"40",x"06",x"00",x"CB",x"47",x"28",x"02",x"CB", -- 0x0F10
    x"C8",x"3A",x"10",x"40",x"CB",x"47",x"28",x"02", -- 0x0F18
    x"CB",x"C0",x"78",x"18",x"C8",x"3A",x"06",x"40", -- 0x0F20
    x"0F",x"30",x"1E",x"3A",x"0D",x"40",x"0F",x"38", -- 0x0F28
    x"26",x"3A",x"10",x"40",x"07",x"07",x"07",x"30", -- 0x0F30
    x"0E",x"DD",x"7E",x"04",x"3C",x"FE",x"D0",x"D0", -- 0x0F38
    x"DD",x"77",x"04",x"DD",x"34",x"24",x"C9",x"07", -- 0x0F40
    x"D0",x"DD",x"7E",x"04",x"3D",x"FE",x"80",x"D8", -- 0x0F48
    x"DD",x"77",x"04",x"DD",x"35",x"24",x"C9",x"3A", -- 0x0F50
    x"11",x"40",x"18",x"D8",x"DD",x"21",x"A0",x"43", -- 0x0F58
    x"CD",x"63",x"1B",x"DD",x"21",x"80",x"43",x"CD", -- 0x0F60
    x"63",x"1B",x"DD",x"34",x"03",x"DD",x"34",x"23", -- 0x0F68
    x"DD",x"7E",x"03",x"FE",x"F0",x"D8",x"DD",x"36", -- 0x0F70
    x"00",x"00",x"DD",x"36",x"01",x"01",x"DD",x"36", -- 0x0F78
    x"02",x"06",x"DD",x"36",x"20",x"00",x"DD",x"36", -- 0x0F80
    x"21",x"01",x"DD",x"36",x"22",x"06",x"C9",x"C9", -- 0x0F88
    x"C9",x"C9",x"21",x"06",x"20",x"22",x"8C",x"43", -- 0x0F90
    x"DD",x"36",x"0E",x"00",x"DD",x"36",x"0F",x"6F", -- 0x0F98
    x"21",x"1E",x"20",x"22",x"AC",x"43",x"DD",x"36", -- 0x0FA0
    x"2E",x"00",x"DD",x"34",x"02",x"3A",x"5F",x"42", -- 0x0FA8
    x"E6",x"03",x"CC",x"DC",x"1F",x"DD",x"21",x"A0", -- 0x0FB0
    x"43",x"CD",x"63",x"1B",x"DD",x"21",x"80",x"43", -- 0x0FB8
    x"CD",x"63",x"1B",x"3A",x"15",x"41",x"A7",x"20", -- 0x0FC0
    x"06",x"DD",x"34",x"04",x"DD",x"34",x"24",x"DD", -- 0x0FC8
    x"35",x"0F",x"C0",x"DD",x"36",x"01",x"00",x"DD", -- 0x0FD0
    x"36",x"21",x"00",x"C9",x"3A",x"17",x"41",x"3C", -- 0x0FD8
    x"E6",x"07",x"32",x"17",x"41",x"C9",x"C9",x"C9", -- 0x0FE0
    x"06",x"28",x"05",x"06",x"2A",x"05",x"06",x"2C", -- 0x0FE8
    x"05",x"06",x"2E",x"05",x"FF",x"E8",x"1F",x"00", -- 0x0FF0
    x"27",x"05",x"00",x"29",x"05",x"00",x"2B",x"05"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
