library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library work;
use work.pace_pkg.all;
use work.video_controller_pkg.all;
use work.sprite_pkg.all;
use work.project_pkg.all;
use work.platform_pkg.all;

entity platform is
  generic
  (
    NUM_INPUT_BYTES   : integer
  );
  port
  (
    -- clocking and reset
    clk_i           : in std_logic_vector(0 to 3);
    reset_i         : in std_logic;

    -- misc I/O
    buttons_i       : in from_BUTTONS_t;
    switches_i      : in from_SWITCHES_t;
    leds_o          : out to_LEDS_t;

    -- controller inputs
    inputs_i        : in from_MAPPED_INPUTS_t(0 to NUM_INPUT_BYTES-1);

    -- FLASH/SRAM
    flash_i         : in from_FLASH_t;
    flash_o         : out to_FLASH_t;
		sram_i					: in from_SRAM_t;
		sram_o					: out to_SRAM_t;

    -- graphics
    
    bitmap_i        : in from_BITMAP_CTL_t;
    bitmap_o        : out to_BITMAP_CTL_t;
    
    tilemap_i       : in from_TILEMAP_CTL_t;
    tilemap_o       : out to_TILEMAP_CTL_t;

    sprite_reg_o    : out to_SPRITE_REG_t;
    sprite_i        : in from_SPRITE_CTL_t;
    sprite_o        : out to_SPRITE_CTL_t;
		spr0_hit				: in std_logic;

    -- various graphics information
    graphics_i      : in from_GRAPHICS_t;
    graphics_o      : out to_GRAPHICS_t;
    
    -- OSD
    osd_i           : in from_OSD_t;
    osd_o           : out to_OSD_t;

    -- sound
    snd_i           : in from_SOUND_t;
    snd_o           : out to_SOUND_t;
    
    -- SPI (flash)
    spi_i           : in from_SPI_t;
    spi_o           : out to_SPI_t;

    -- serial
    ser_i           : in from_SERIAL_t;
    ser_o           : out to_SERIAL_t;

    -- general purpose I/O
    gp_i            : in from_GP_t;
    gp_o            : out to_GP_t
  );

end platform;

architecture SYN of platform is

	alias clk_30M					: std_logic is clk_i(0);
	alias clk_video 			: std_logic is clk_i(1);
	
	signal reset_n				: std_logic;
	
  -- uP signals  
  signal clk_1M5_ena		: std_logic;
  signal up_addr        : std_logic_vector(23 downto 0);
	alias addr_bus				: std_logic_vector(13 downto 0) is up_addr(13 downto 0);
  signal up_datai       : std_logic_vector(7 downto 0);
  signal up_datao       : std_logic_vector(7 downto 0);
  signal up_rw_n				: std_logic;
  signal up_irq_n				: std_logic;
	                        
  -- ROM signals        
	signal rom_cs					: std_logic;
  signal rom_data      	: std_logic_vector(7 downto 0);
                        
  -- keyboard signals
	                        
  -- VRAM signals       
	signal vram_cs				: std_logic;
	signal vram_wr				: std_logic;
	signal vram_addr			: std_logic_vector(9 downto 0);
  signal vram_datao     : std_logic_vector(7 downto 0);
                        
  -- RAM signals        
  signal wram_cs        : std_logic;
	signal wram_wr				: std_logic;
  alias wram_datao     	: std_logic_vector(7 downto 0) is sram_i.d(7 downto 0);

  -- RAM signals        
  signal cram_cs        : std_logic;
  signal cram_wr        : std_logic;
	signal cram0_wr				: std_logic;
	signal cram1_wr				: std_logic;
	signal cram0_datao		: std_logic_vector(7 downto 0);
	signal cram1_datao		: std_logic_vector(7 downto 0);
	
  -- other signals      
  signal dip_cs 				: std_logic;
  signal in0_cs 				: std_logic;
  signal in1_cs 				: std_logic;
  signal in2_cs 				: std_logic;
  signal in3_cs 				: std_logic;
	signal pokey_cs 			: std_logic;
	signal sprite_cs      : std_logic;
  signal intack_wr			: std_logic;
	signal vblank_n				: std_logic;			-- should be vsync, but we don't have that
	signal vblank_fake		: std_logic;			-- generated by intgen, not video controller
	
	signal newtileAddr		: std_logic_vector(11 downto 0);
	
begin

	reset_n <= not reset_i;
	vblank_n <= not graphics_i.vblank;
	
  -- centipede A15 & A14 aren't connected on the PCB
  -- chip select logic

	-- WRAM $0000-$03FF
	-- SPRITE_RAM $07C0-$07FF (use SRAM atm)
	-- atari_vg_earom $1700-$173F
	wram_cs <= 	'1' when STD_MATCH(addr_bus, "0000----------") else 
							'1' when STD_MATCH(addr_bus, "00011111------") else
							'1' when STD_MATCH(addr_bus, "01011100------") else
							'0';
	-- VRAM $0400-$07BF
	vram_cs <= 	'1' when addr_bus(13 downto 10) = "0001" and addr_bus(9 downto 6) /= "1111" else '0';
	-- DIP0 $0800
  dip_cs <= 	'1' when STD_MATCH(addr_bus, "00100000000000") else '0';
	-- IN0 $0C00 (analog?)
  in0_cs <= 	'1' when STD_MATCH(addr_bus, "00110000000000") else '0';
	-- IN1 $0C01 (digital)
  in1_cs <= 	'1' when STD_MATCH(addr_bus, "00110000000001") else '0';
	-- IN2 $0C02 (analog?)
  in2_cs <= 	'1' when STD_MATCH(addr_bus, "00110000000010") else '0';
	-- IN3 $0C03 (digital)
  in3_cs <= 	'1' when STD_MATCH(addr_bus, "00110000000011") else '0';
	-- POKEY $1000-$100F
	pokey_cs <=	'1' when STD_MATCH(addr_bus, "0100000000----") else '0';
	-- ROM $2000-$3FFF
  rom_cs <= 	'1' when STD_MATCH(addr_bus, "1-------------") else '0';

	-- memory read mux
	uP_datai <= vram_datao when vram_cs = '1' else
							not switches_i(7 downto 0) when dip_cs = '1' else
							(inputs_i(0).d(7) & vblank_fake & inputs_i(0).d(5 downto 0)) when in0_cs = '1' else
							inputs_i(1).d when in1_cs = '1' else
							inputs_i(2).d when in2_cs = '1' else
							X"00" when in3_cs = '1' else
							snd_i.d when pokey_cs = '1' else
							rom_data when rom_cs = '1' else
							wram_datao;

  snd_o.rd <= up_rw_n and pokey_cs;

	-- wram $0000-$03FF
	-- sprite_wr $07C0-$07FF
	-- atari_vg_earom $1600-$163F
  -- atari_vg_earom_ctrl $1680
	-- * handled below
  -- vram_wr $0400-$07BF
	vram_wr <= not up_rw_n and vram_cs;
	-- sprite_wr $07C0-$07FF
  sprite_cs <= '1' when addr_bus(13 downto 6) = "00011111" else '0';
	-- POKEY $1000-$100F
  snd_o.wr <= not up_rw_n and pokey_cs;
	-- palette ram $1400-$140F
  cram_wr <= not up_rw_n when addr_bus(13 downto 4) = "0101000000" else '0';
	-- intack_wr $1800
  intack_wr <= not up_rw_n when addr_bus = "01100000000000" else '0';

  snd_o.a <= addr_bus(snd_o.a'range);
  snd_o.d <= up_datao;

  -- sprite register address
  -- sprite registers for sprite #0 @ $00,$10,$20,$30
  -- sprite registers for sprite #1 @ $01,$11,$21,$31
  sprite_reg_o.clk <= clk_30M;
  sprite_reg_o.clk_ena <= clk_1M5_ena;
  sprite_reg_o.a <= addr_bus(7 downto 6) & addr_bus(3 downto 0) & addr_bus(5 downto 4);
  sprite_reg_o.d <= up_datao;
  sprite_reg_o.wr <= not up_rw_n and sprite_cs;
  
	-- mangle sprite address according to tile layout
	newTileAddr <=  tilemap_i.tile_a(11 downto 5) & tilemap_i.tile_a(3 downto 1) & 
                  tilemap_i.tile_a(4) & tilemap_i.tile_a(0);

  -- SRAM signals (may or may not be used)
  sram_o.a <= std_logic_vector(resize(unsigned(addr_bus), sram_o.a'length));
  sram_o.d <= std_logic_vector(resize(unsigned(up_datao), sram_o.d'length));
	sram_o.be <= std_logic_vector(to_unsigned(1, sram_o.be'length));
  sram_o.cs <= '1';
  sram_o.oe <= wram_cs and up_rw_n;
  sram_o.we <= wram_cs and not up_rw_n;
	
  -- unused outputs
  flash_o <= NULL_TO_FLASH;
  bitmap_o <= NULL_TO_BITMAP_CTL;
  graphics_o <= NULL_TO_GRAPHICS;
  spi_o <= NULL_TO_SPI;
  ser_o <= NULL_TO_SERIAL;
  osd_o <= NULL_TO_OSD;
	leds_o <= std_logic_vector(resize(unsigned(inputs_i(0).d), leds_o'length));
	gp_o <= (others => '0');
	
  --
  -- COMPONENT INSTANTIATION
  --

	-- generate CPU clock enable (1M5Hz from 30MHz)
	clk_en_inst : entity work.clk_div
		generic map
		(
			DIVISOR		=> 20
		)
		port map
		(
			clk				=> clk_30M,
			reset			=> reset_i,
			clk_en		=> clk_1M5_ena
		);

	up_inst : entity work.T65
		port map
		(
			Mode    		=> "00",	-- 6502
			Res_n   		=> reset_n,
			Enable  		=> clk_1M5_ena,
			Clk     		=> clk_30M,
			Rdy     		=> '1',
			Abort_n 		=> '1',
			IRQ_n   		=> up_irq_n,
			NMI_n   		=> '1',
			SO_n    		=> '1',
			R_W_n   		=> up_rw_n,
			Sync    		=> open,
			EF      		=> open,
			MF      		=> open,
			XF      		=> open,
			ML_n    		=> open,
			VP_n    		=> open,
			VDA     		=> open,
			VPA     		=> open,
			A       		=> up_addr,
			DI      		=> up_datai,
			DO      		=> up_datao
		);

	rom_inst : entity work.sprom
		generic map
		(
			init_file		=> "../../../../src/platform/centiped/roms/rom0.hex",
			numwords_a	=> 8192,
			widthad_a		=> 13
		)
		port map
		(
			clock			=> clk_30M,
			address		=> addr_bus(12 downto 0),
			q					=> rom_data
		);
	
	vram_inst : entity work.dpram
		-- wren_a *MUST* be GND for CYCLONEII_SAFE_WRITE=VERIFIED_SAFE
		generic map
		(
			init_file		=> "../../../../src/platform/centiped/roms/vram.hex",
			numwords_a	=> 1024,
			widthad_a		=> 10
		)
		port map
		(
			clock_b			=> clk_30M,
			address_b		=> addr_bus(9 downto 0),
			wren_b			=> vram_wr,
			data_b			=> up_datao,
			q_b					=> vram_datao,

			clock_a			=> clk_video,
			address_a		=> vram_addr,
			wren_a			=> '0',
			data_a			=> (others => 'X'),
			q_a					=> tilemap_o.map_d(7 downto 0)
		);
	tilemap_o.map_d(15 downto 8) <= (others => '0');
	
	vrammapper_inst : entity work.vramMapper
		port map
		(
	    clk     => clk_video,

	    inAddr  => tilemap_i.map_a(12 downto 0),
	    outAddr => vram_addr
		);

	cram0_wr <= cram_wr and not addr_bus(0);
	
	-- wren_a *MUST* be GND for CYCLONEII_SAFE_WRITE=VERIFIED_SAFE
	cram_inst_0 : entity work.dpram
		generic map
		(
			numwords_a			=> 128,
			widthad_a				=> 7
		)
		port map
		(
			clock_b					=> clk_30M,
			address_b				=> addr_bus(7 downto 1),
			wren_b					=> cram0_wr,
			data_b					=> up_datao,
			q_b							=> cram0_datao,
			
			clock_a					=> clk_video,
			address_a				=> tilemap_i.attr_a(7 downto 1),
			wren_a					=> '0',
			data_a					=> (others => 'X'),
			q_a							=> tilemap_o.attr_d(7 downto 0)
		);

	cram1_wr <= cram_wr and addr_bus(0);

	-- wren_a *MUST* be GND for CYCLONEII_SAFE_WRITE=VERIFIED_SAFE
	cram_inst_1 : entity work.dpram
		generic map
		(
			numwords_a			=> 128,
			widthad_a				=> 7
		)
		port map
		(
			clock_b					=> clk_30M,
			address_b				=> addr_bus(7 downto 1),
			wren_b					=> cram1_wr,
			data_b					=> up_datao,
			q_b							=> cram1_datao,
			
			clock_a					=> clk_video,
			address_a				=> tilemap_i.attr_a(7 downto 1),
			wren_a					=> '0',
			data_a					=> (others => 'X'),
			q_a							=> tilemap_o.attr_d(15 downto 8)
		);

	intgen_inst : entity work.intGen
		port map
		(
	    clk       	=> clk_30M,
	    reset     	=> reset_i,

	    -- inputs
	    vsync_n   	=> vblank_n,
	    intack    	=> intack_wr,

	    -- outputs
	    vblank    	=> vblank_fake,
	    irq_n     	=> up_irq_n
		);

	gfxrom_inst : entity work.dprom_2r
		generic map
		(
			init_file		=> "../../../../src/platform/centiped/roms/gfxrom.hex",
			numwords_a	=> 4096,
			widthad_a		=> 12,
			numwords_b	=> 1024,
			widthad_b		=> 10,
			width_b			=> 32
		)
		port map
		(
			clock										=> clk_video,
			address_a								=> newtileaddr(11 downto 0),
			q_a											=> tilemap_o.tile_d,
			
			address_b								=> sprite_i.a(9 downto 0),
			q_b(31 downto 24)				=> sprite_o.d(7 downto 0),
			q_b(23 downto 16)				=> sprite_o.d(15 downto 8),
			q_b(15 downto 8)				=> sprite_o.d(23 downto 16),
			q_b(7 downto 0)					=> sprite_o.d(31 downto 24)
		);

end SYN;
