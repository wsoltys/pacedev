-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_PGM_23 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_PGM_23 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"15",x"14",x"19",x"24",x"24",x"19",x"1D",x"15", -- 0x0000
    x"10",x"10",x"20",x"15",x"22",x"20",x"25",x"23", -- 0x0008
    x"18",x"10",x"23",x"24",x"11",x"22",x"24",x"10", -- 0x0010
    x"12",x"25",x"24",x"24",x"1F",x"1E",x"1F",x"1E", -- 0x0018
    x"15",x"10",x"1F",x"22",x"10",x"24",x"27",x"1F", -- 0x0020
    x"10",x"20",x"1C",x"11",x"29",x"15",x"22",x"10", -- 0x0028
    x"1F",x"1E",x"1C",x"29",x"12",x"1F",x"1E",x"25", -- 0x0030
    x"23",x"10",x"15",x"28",x"24",x"22",x"11",x"10", -- 0x0038
    x"16",x"22",x"1F",x"17",x"23",x"10",x"11",x"16", -- 0x0040
    x"24",x"15",x"22",x"10",x"20",x"24",x"23",x"FF", -- 0x0048
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0060
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0068
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0070
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0078
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0080
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0088
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0090
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0098
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0100
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0108
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0110
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0118
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0120
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0128
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0130
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0138
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0140
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0148
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0150
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0158
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0160
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0168
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0170
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0178
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0180
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0188
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0190
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0198
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0200
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0208
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0210
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0218
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0220
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0228
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0230
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0238
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0240
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0248
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0250
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0258
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0260
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0268
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0270
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0278
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0280
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0288
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0290
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0298
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0300
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0308
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0310
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0318
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0320
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0328
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0330
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0338
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0340
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0348
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0350
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0358
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0360
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0368
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0370
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0378
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0380
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0388
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0390
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0398
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0400
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0408
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0410
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0418
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0420
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0428
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0430
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0438
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0440
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0448
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0450
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0458
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0460
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0468
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0470
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0478
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0480
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0488
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0490
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0498
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0500
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0508
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0510
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0518
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0520
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0528
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0530
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0538
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0540
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0548
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0550
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0558
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0560
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0568
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0570
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0578
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0580
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0588
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0590
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0598
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0600
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0608
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0610
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0618
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0620
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0628
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0630
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0638
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0640
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0648
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0650
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0658
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0660
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0668
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0670
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0678
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0680
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0688
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0690
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0698
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0700
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0708
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0710
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0718
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0720
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0728
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0730
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0738
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F8
    x"3A",x"86",x"83",x"A7",x"C2",x"B0",x"19",x"21", -- 0x0800
    x"D8",x"83",x"7E",x"B7",x"C0",x"36",x"80",x"2D", -- 0x0808
    x"7E",x"34",x"21",x"1F",x"18",x"07",x"4F",x"06", -- 0x0810
    x"00",x"09",x"46",x"23",x"66",x"68",x"E9",x"3B", -- 0x0818
    x"18",x"68",x"18",x"7A",x"18",x"97",x"18",x"B4", -- 0x0820
    x"18",x"D7",x"18",x"DD",x"18",x"21",x"19",x"38", -- 0x0828
    x"19",x"49",x"19",x"5A",x"19",x"77",x"19",x"88", -- 0x0830
    x"19",x"A5",x"19",x"3E",x"06",x"32",x"17",x"80", -- 0x0838
    x"32",x"19",x"80",x"32",x"1B",x"80",x"32",x"1D", -- 0x0840
    x"80",x"3E",x"03",x"32",x"21",x"80",x"32",x"23", -- 0x0848
    x"80",x"32",x"25",x"80",x"32",x"27",x"80",x"3E", -- 0x0850
    x"01",x"32",x"2B",x"80",x"32",x"2D",x"80",x"32", -- 0x0858
    x"31",x"80",x"32",x"2F",x"80",x"C3",x"15",x"19", -- 0x0860
    x"11",x"B5",x"19",x"06",x"18",x"21",x"88",x"AB", -- 0x0868
    x"EF",x"06",x"1B",x"21",x"89",x"AB",x"EF",x"C3", -- 0x0870
    x"15",x"19",x"11",x"E8",x"19",x"06",x"14",x"21", -- 0x0878
    x"8B",x"AB",x"EF",x"06",x"1A",x"21",x"8C",x"AB", -- 0x0880
    x"EF",x"06",x"15",x"21",x"8D",x"AB",x"EF",x"06", -- 0x0888
    x"1A",x"21",x"8E",x"AB",x"EF",x"18",x"7E",x"11", -- 0x0890
    x"45",x"1A",x"06",x"16",x"21",x"90",x"AB",x"EF", -- 0x0898
    x"06",x"15",x"21",x"91",x"AB",x"EF",x"06",x"14", -- 0x08A0
    x"21",x"92",x"AB",x"EF",x"06",x"0A",x"21",x"93", -- 0x08A8
    x"AB",x"EF",x"18",x"61",x"11",x"8E",x"1A",x"06", -- 0x08B0
    x"15",x"21",x"95",x"AB",x"EF",x"06",x"19",x"21", -- 0x08B8
    x"96",x"AB",x"EF",x"06",x"14",x"21",x"97",x"AB", -- 0x08C0
    x"EF",x"06",x"0E",x"21",x"98",x"AB",x"EF",x"3E", -- 0x08C8
    x"A0",x"32",x"86",x"83",x"C3",x"1B",x"19",x"21", -- 0x08D0
    x"D8",x"83",x"36",x"C0",x"C9",x"CD",x"79",x"07", -- 0x08D8
    x"3E",x"06",x"32",x"0F",x"80",x"32",x"15",x"80", -- 0x08E0
    x"32",x"1B",x"80",x"32",x"25",x"80",x"32",x"2B", -- 0x08E8
    x"80",x"32",x"33",x"80",x"3E",x"03",x"32",x"0D", -- 0x08F0
    x"80",x"32",x"13",x"80",x"32",x"19",x"80",x"32", -- 0x08F8
    x"21",x"80",x"32",x"23",x"80",x"32",x"29",x"80", -- 0x0900
    x"32",x"2F",x"80",x"32",x"31",x"80",x"AF",x"32", -- 0x0908
    x"0B",x"80",x"32",x"1F",x"80",x"21",x"D8",x"83", -- 0x0910
    x"36",x"80",x"C9",x"21",x"D8",x"83",x"36",x"F0", -- 0x0918
    x"C9",x"11",x"DE",x"1A",x"06",x"12",x"21",x"85", -- 0x0920
    x"AB",x"EF",x"06",x"13",x"21",x"86",x"AB",x"EF", -- 0x0928
    x"06",x"0B",x"21",x"87",x"AB",x"EF",x"18",x"DD", -- 0x0930
    x"11",x"0E",x"1B",x"06",x"15",x"21",x"89",x"AB", -- 0x0938
    x"EF",x"06",x"0B",x"21",x"8A",x"AB",x"EF",x"18", -- 0x0940
    x"CC",x"11",x"2E",x"1B",x"06",x"1A",x"21",x"8C", -- 0x0948
    x"AB",x"EF",x"06",x"1A",x"21",x"8D",x"AB",x"EF", -- 0x0950
    x"18",x"BB",x"11",x"62",x"1B",x"06",x"18",x"21", -- 0x0958
    x"8F",x"AB",x"EF",x"06",x"12",x"21",x"90",x"AB", -- 0x0960
    x"EF",x"06",x"0C",x"21",x"91",x"AB",x"EF",x"06", -- 0x0968
    x"0C",x"21",x"92",x"AB",x"EF",x"18",x"9E",x"11", -- 0x0970
    x"A4",x"1B",x"06",x"13",x"21",x"94",x"AB",x"EF", -- 0x0978
    x"06",x"0C",x"21",x"95",x"AB",x"EF",x"18",x"8D", -- 0x0980
    x"11",x"C3",x"1B",x"06",x"13",x"21",x"97",x"AB", -- 0x0988
    x"EF",x"06",x"14",x"21",x"98",x"AB",x"EF",x"06", -- 0x0990
    x"0D",x"21",x"99",x"AB",x"EF",x"3E",x"A0",x"32", -- 0x0998
    x"86",x"83",x"C3",x"1B",x"19",x"3E",x"03",x"32", -- 0x09A0
    x"D6",x"83",x"21",x"D8",x"83",x"36",x"C0",x"C9", -- 0x09A8
    x"21",x"86",x"83",x"35",x"C9",x"1D",x"1F",x"26", -- 0x09B0
    x"15",x"10",x"16",x"22",x"1F",x"17",x"10",x"26", -- 0x09B8
    x"15",x"22",x"24",x"19",x"13",x"11",x"1C",x"1C", -- 0x09C0
    x"29",x"10",x"1F",x"22",x"10",x"18",x"1F",x"22", -- 0x09C8
    x"19",x"2A",x"1F",x"1E",x"24",x"11",x"1C",x"1C", -- 0x09D0
    x"29",x"10",x"25",x"23",x"19",x"1E",x"17",x"10", -- 0x09D8
    x"1A",x"1F",x"29",x"23",x"24",x"19",x"13",x"1B", -- 0x09E0
    x"1F",x"12",x"1A",x"15",x"13",x"24",x"10",x"19", -- 0x09E8
    x"23",x"10",x"24",x"1F",x"10",x"23",x"11",x"16", -- 0x09F0
    x"15",x"1C",x"29",x"10",x"1D",x"11",x"1E",x"15", -- 0x09F8
    x"25",x"26",x"15",x"22",x"10",x"16",x"22",x"1F", -- 0x0A00
    x"17",x"10",x"24",x"1F",x"10",x"19",x"24",x"23", -- 0x0A08
    x"10",x"18",x"1F",x"1D",x"15",x"10",x"27",x"19", -- 0x0A10
    x"24",x"18",x"19",x"1E",x"10",x"11",x"1C",x"1C", -- 0x0A18
    x"1F",x"24",x"24",x"15",x"14",x"10",x"24",x"19", -- 0x0A20
    x"1D",x"15",x"10",x"2B",x"23",x"19",x"28",x"24", -- 0x0A28
    x"29",x"10",x"12",x"15",x"11",x"24",x"23",x"10", -- 0x0A30
    x"1F",x"1E",x"10",x"24",x"18",x"15",x"10",x"24", -- 0x0A38
    x"19",x"1D",x"15",x"22",x"2B",x"13",x"22",x"1F", -- 0x0A40
    x"23",x"23",x"10",x"18",x"19",x"17",x"18",x"27", -- 0x0A48
    x"11",x"29",x"10",x"27",x"19",x"24",x"18",x"1F", -- 0x0A50
    x"25",x"24",x"10",x"17",x"15",x"24",x"24",x"19", -- 0x0A58
    x"1E",x"17",x"10",x"22",x"25",x"1E",x"10",x"1F", -- 0x0A60
    x"26",x"15",x"22",x"10",x"11",x"1E",x"14",x"10", -- 0x0A68
    x"13",x"22",x"1F",x"23",x"23",x"10",x"22",x"19", -- 0x0A70
    x"26",x"15",x"22",x"10",x"27",x"19",x"24",x"18", -- 0x0A78
    x"1F",x"25",x"24",x"10",x"16",x"11",x"1C",x"1C", -- 0x0A80
    x"19",x"1E",x"17",x"10",x"19",x"1E",x"11",x"26", -- 0x0A88
    x"1F",x"19",x"14",x"10",x"24",x"22",x"11",x"16", -- 0x0A90
    x"16",x"19",x"13",x"10",x"14",x"15",x"11",x"14", -- 0x0A98
    x"1C",x"29",x"10",x"23",x"1E",x"11",x"1B",x"15", -- 0x0AA0
    x"23",x"10",x"1F",x"24",x"24",x"15",x"22",x"23", -- 0x0AA8
    x"10",x"13",x"22",x"1F",x"13",x"1F",x"14",x"19", -- 0x0AB0
    x"1C",x"15",x"23",x"10",x"11",x"1E",x"14",x"10", -- 0x0AB8
    x"24",x"18",x"15",x"10",x"24",x"22",x"15",x"11", -- 0x0AC0
    x"13",x"18",x"15",x"22",x"1F",x"25",x"23",x"10", -- 0x0AC8
    x"14",x"19",x"26",x"19",x"1E",x"17",x"10",x"24", -- 0x0AD0
    x"25",x"22",x"24",x"1C",x"15",x"23",x"20",x"1F", -- 0x0AD8
    x"19",x"1E",x"24",x"23",x"10",x"11",x"22",x"15", -- 0x0AE0
    x"10",x"23",x"13",x"1F",x"22",x"15",x"14",x"10", -- 0x0AE8
    x"16",x"1F",x"22",x"10",x"15",x"11",x"13",x"18", -- 0x0AF0
    x"10",x"23",x"11",x"16",x"15",x"10",x"1A",x"25", -- 0x0AF8
    x"1D",x"20",x"10",x"2B",x"01",x"00",x"10",x"20", -- 0x0B00
    x"1F",x"19",x"1E",x"24",x"23",x"2B",x"23",x"11", -- 0x0B08
    x"16",x"15",x"1C",x"29",x"10",x"11",x"22",x"22", -- 0x0B10
    x"19",x"26",x"19",x"1E",x"17",x"10",x"18",x"1F", -- 0x0B18
    x"1D",x"15",x"10",x"2B",x"05",x"00",x"10",x"20", -- 0x0B20
    x"1F",x"19",x"1E",x"24",x"23",x"2B",x"11",x"1E", -- 0x0B28
    x"14",x"10",x"16",x"1F",x"22",x"10",x"12",x"15", -- 0x0B30
    x"11",x"24",x"19",x"1E",x"17",x"10",x"24",x"18", -- 0x0B38
    x"15",x"10",x"24",x"19",x"1D",x"15",x"22",x"10", -- 0x0B40
    x"2B",x"01",x"00",x"10",x"20",x"1F",x"19",x"1E", -- 0x0B48
    x"24",x"23",x"10",x"20",x"15",x"22",x"10",x"12", -- 0x0B50
    x"15",x"11",x"24",x"10",x"23",x"11",x"26",x"15", -- 0x0B58
    x"14",x"2B",x"12",x"1F",x"1E",x"25",x"23",x"10", -- 0x0B60
    x"20",x"1F",x"19",x"1E",x"24",x"23",x"10",x"11", -- 0x0B68
    x"22",x"15",x"10",x"23",x"13",x"1F",x"22",x"15", -- 0x0B70
    x"14",x"10",x"12",x"29",x"10",x"15",x"23",x"13", -- 0x0B78
    x"1F",x"22",x"24",x"19",x"1E",x"17",x"10",x"18", -- 0x0B80
    x"1F",x"1D",x"15",x"10",x"11",x"10",x"1C",x"11", -- 0x0B88
    x"14",x"29",x"10",x"16",x"22",x"1F",x"17",x"10", -- 0x0B90
    x"2B",x"02",x"00",x"00",x"10",x"20",x"1F",x"19", -- 0x0B98
    x"1E",x"24",x"23",x"2B",x"17",x"1F",x"12",x"12", -- 0x0BA0
    x"1C",x"19",x"1E",x"17",x"10",x"11",x"1E",x"10", -- 0x0BA8
    x"19",x"1E",x"23",x"15",x"13",x"24",x"10",x"2B", -- 0x0BB0
    x"02",x"00",x"00",x"10",x"20",x"1F",x"19",x"1E", -- 0x0BB8
    x"24",x"23",x"2B",x"11",x"1E",x"14",x"10",x"23", -- 0x0BC0
    x"11",x"16",x"15",x"1C",x"29",x"10",x"17",x"15", -- 0x0BC8
    x"24",x"24",x"19",x"1E",x"17",x"10",x"11",x"1C", -- 0x0BD0
    x"1C",x"10",x"16",x"19",x"26",x"15",x"10",x"16", -- 0x0BD8
    x"22",x"1F",x"17",x"23",x"10",x"18",x"1F",x"1D", -- 0x0BE0
    x"15",x"10",x"2B",x"01",x"00",x"00",x"00",x"10", -- 0x0BE8
    x"20",x"1F",x"19",x"1E",x"24",x"23",x"2B",x"FF", -- 0x0BF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF8
    x"3A",x"B7",x"83",x"FE",x"03",x"38",x"2A",x"3A", -- 0x0C00
    x"FD",x"83",x"3D",x"20",x"06",x"DD",x"21",x"40", -- 0x0C08
    x"84",x"18",x"04",x"DD",x"21",x"60",x"84",x"FD", -- 0x0C10
    x"21",x"48",x"80",x"CD",x"49",x"1C",x"3A",x"B7", -- 0x0C18
    x"83",x"FE",x"06",x"38",x"07",x"11",x"10",x"00", -- 0x0C20
    x"DD",x"19",x"FD",x"21",x"50",x"80",x"CD",x"49", -- 0x0C28
    x"1C",x"3A",x"FD",x"83",x"3D",x"20",x"06",x"DD", -- 0x0C30
    x"21",x"80",x"84",x"18",x"04",x"DD",x"21",x"90", -- 0x0C38
    x"84",x"FD",x"21",x"58",x"80",x"CD",x"13",x"1E", -- 0x0C40
    x"C9",x"CD",x"FA",x"1C",x"CD",x"59",x"1C",x"CD", -- 0x0C48
    x"89",x"1C",x"CD",x"83",x"1D",x"CD",x"E8",x"1D", -- 0x0C50
    x"C9",x"DD",x"35",x"08",x"C0",x"DD",x"36",x"08", -- 0x0C58
    x"0C",x"DD",x"7E",x"06",x"B7",x"C8",x"3D",x"20", -- 0x0C60
    x"02",x"3E",x"04",x"DD",x"77",x"06",x"6F",x"26", -- 0x0C68
    x"00",x"11",x"65",x"1F",x"19",x"7E",x"DD",x"B6", -- 0x0C70
    x"05",x"FD",x"77",x"01",x"3C",x"FD",x"77",x"05", -- 0x0C78
    x"FD",x"36",x"02",x"04",x"FD",x"36",x"06",x"04", -- 0x0C80
    x"C9",x"DD",x"7E",x"06",x"B7",x"C8",x"3A",x"2C", -- 0x0C88
    x"84",x"B7",x"C0",x"DD",x"35",x"09",x"C0",x"DD", -- 0x0C90
    x"36",x"09",x"08",x"FD",x"7E",x"03",x"FE",x"60", -- 0x0C98
    x"30",x"2A",x"DD",x"36",x"07",x"01",x"DD",x"7E", -- 0x0CA0
    x"05",x"B7",x"C2",x"BD",x"1C",x"3A",x"14",x"80", -- 0x0CA8
    x"DD",x"96",x"00",x"D8",x"FD",x"BE",x"00",x"30", -- 0x0CB0
    x"2A",x"DD",x"34",x"02",x"C9",x"3A",x"14",x"80", -- 0x0CB8
    x"DD",x"96",x"01",x"FD",x"BE",x"00",x"38",x"1B", -- 0x0CC0
    x"DD",x"35",x"02",x"C9",x"DD",x"36",x"07",x"01", -- 0x0CC8
    x"DD",x"7E",x"05",x"B7",x"28",x"04",x"3E",x"02", -- 0x0CD0
    x"18",x"02",x"3E",x"FE",x"DD",x"86",x"03",x"DD", -- 0x0CD8
    x"77",x"03",x"C9",x"DD",x"7E",x"05",x"EE",x"80", -- 0x0CE0
    x"DD",x"77",x"05",x"FD",x"7E",x"04",x"FD",x"77", -- 0x0CE8
    x"00",x"FD",x"7E",x"01",x"EE",x"80",x"FD",x"77", -- 0x0CF0
    x"01",x"C9",x"3A",x"B7",x"83",x"FE",x"03",x"D8", -- 0x0CF8
    x"4F",x"DD",x"35",x"0A",x"C0",x"DD",x"7E",x"06", -- 0x0D00
    x"B7",x"C0",x"CD",x"11",x"0B",x"47",x"79",x"87", -- 0x0D08
    x"87",x"87",x"C6",x"80",x"B8",x"D8",x"CD",x"11", -- 0x0D10
    x"0B",x"E6",x"03",x"28",x"1D",x"0E",x"40",x"21", -- 0x0D18
    x"76",x"82",x"7E",x"0F",x"0F",x"C6",x"24",x"57", -- 0x0D20
    x"2C",x"2C",x"46",x"3A",x"14",x"80",x"D6",x"10", -- 0x0D28
    x"38",x"08",x"91",x"38",x"19",x"92",x"38",x"02", -- 0x0D30
    x"10",x"F8",x"DD",x"36",x"04",x"7E",x"CD",x"11", -- 0x0D38
    x"0B",x"0F",x"38",x"1E",x"DD",x"36",x"05",x"00", -- 0x0D40
    x"DD",x"36",x"03",x"F0",x"18",x"1C",x"81",x"47", -- 0x0D48
    x"3A",x"14",x"80",x"DD",x"77",x"02",x"90",x"DD", -- 0x0D50
    x"77",x"01",x"81",x"DD",x"77",x"00",x"DD",x"36", -- 0x0D58
    x"04",x"4E",x"DD",x"36",x"05",x"80",x"DD",x"36", -- 0x0D60
    x"03",x"00",x"DD",x"36",x"06",x"01",x"DD",x"36", -- 0x0D68
    x"08",x"0B",x"DD",x"36",x"09",x"08",x"3A",x"71", -- 0x0D70
    x"83",x"B7",x"C0",x"3C",x"32",x"71",x"83",x"3E", -- 0x0D78
    x"90",x"DF",x"C9",x"DD",x"7E",x"06",x"B7",x"C8", -- 0x0D80
    x"CD",x"76",x"1D",x"DD",x"7E",x"04",x"FE",x"60", -- 0x0D88
    x"30",x"0C",x"3A",x"14",x"80",x"DD",x"96",x"02", -- 0x0D90
    x"4F",x"FD",x"77",x"00",x"18",x"06",x"DD",x"4E", -- 0x0D98
    x"03",x"FD",x"71",x"00",x"DD",x"7E",x"04",x"FD", -- 0x0DA0
    x"77",x"03",x"FD",x"77",x"07",x"DD",x"7E",x"05", -- 0x0DA8
    x"B7",x"20",x"0A",x"3E",x"0F",x"81",x"FD",x"77", -- 0x0DB0
    x"04",x"3C",x"C0",x"18",x"09",x"3E",x"F1",x"81", -- 0x0DB8
    x"FD",x"77",x"04",x"79",x"B7",x"C0",x"DD",x"7E", -- 0x0DC0
    x"07",x"B7",x"C8",x"DD",x"E5",x"E1",x"54",x"5D", -- 0x0DC8
    x"1C",x"01",x"0F",x"00",x"70",x"ED",x"B0",x"01", -- 0x0DD0
    x"07",x"00",x"FD",x"E5",x"E1",x"54",x"5D",x"1C", -- 0x0DD8
    x"70",x"ED",x"B0",x"DD",x"36",x"0A",x"20",x"C9", -- 0x0DE0
    x"DD",x"7E",x"06",x"B7",x"C8",x"DD",x"7E",x"04", -- 0x0DE8
    x"C6",x"02",x"21",x"47",x"80",x"BE",x"C0",x"DD", -- 0x0DF0
    x"7E",x"05",x"B7",x"FD",x"7E",x"00",x"21",x"44", -- 0x0DF8
    x"80",x"28",x"02",x"C6",x"10",x"96",x"D8",x"FE", -- 0x0E00
    x"10",x"D0",x"3E",x"01",x"32",x"04",x"80",x"32", -- 0x0E08
    x"2C",x"84",x"C9",x"CD",x"A3",x"1E",x"CD",x"3B", -- 0x0E10
    x"1E",x"CD",x"23",x"1E",x"CD",x"38",x"1F",x"CD", -- 0x0E18
    x"8B",x"1E",x"C9",x"DD",x"7E",x"06",x"B7",x"C8", -- 0x0E20
    x"DD",x"6E",x"0B",x"26",x"80",x"7E",x"DD",x"96", -- 0x0E28
    x"02",x"FD",x"77",x"00",x"DD",x"7E",x"04",x"FD", -- 0x0E30
    x"77",x"03",x"C9",x"DD",x"7E",x"06",x"B7",x"C8", -- 0x0E38
    x"DD",x"35",x"09",x"C0",x"DD",x"36",x"09",x"08", -- 0x0E40
    x"DD",x"6E",x"0B",x"26",x"80",x"DD",x"7E",x"05", -- 0x0E48
    x"B7",x"28",x"0D",x"7E",x"DD",x"96",x"00",x"FD", -- 0x0E50
    x"BE",x"00",x"30",x"11",x"DD",x"34",x"02",x"C9", -- 0x0E58
    x"7E",x"DD",x"96",x"01",x"FD",x"BE",x"00",x"38", -- 0x0E60
    x"04",x"DD",x"35",x"02",x"C9",x"3A",x"04",x"80", -- 0x0E68
    x"B7",x"C0",x"DD",x"E5",x"E1",x"54",x"5D",x"1C", -- 0x0E70
    x"01",x"0F",x"00",x"70",x"ED",x"B0",x"21",x"58", -- 0x0E78
    x"80",x"11",x"59",x"80",x"01",x"03",x"00",x"70", -- 0x0E80
    x"ED",x"B0",x"C9",x"DD",x"7E",x"06",x"B7",x"C8", -- 0x0E88
    x"21",x"69",x"1F",x"4F",x"06",x"00",x"09",x"7E", -- 0x0E90
    x"DD",x"B6",x"05",x"FD",x"77",x"01",x"FD",x"36", -- 0x0E98
    x"02",x"02",x"C9",x"3A",x"B7",x"83",x"FE",x"03", -- 0x0EA0
    x"D8",x"4F",x"DD",x"7E",x"06",x"B7",x"C0",x"CD", -- 0x0EA8
    x"11",x"0B",x"47",x"79",x"87",x"87",x"87",x"C6", -- 0x0EB0
    x"80",x"B8",x"D8",x"0E",x"40",x"CD",x"11",x"0B", -- 0x0EB8
    x"E6",x"07",x"FE",x"05",x"D0",x"4F",x"0F",x"0F", -- 0x0EC0
    x"0F",x"0F",x"C6",x"30",x"DD",x"77",x"04",x"CD", -- 0x0EC8
    x"11",x"0B",x"47",x"79",x"87",x"5F",x"16",x"00", -- 0x0ED0
    x"21",x"76",x"1F",x"19",x"5E",x"2C",x"6E",x"26", -- 0x0ED8
    x"80",x"DD",x"75",x"0B",x"7E",x"57",x"79",x"87", -- 0x0EE0
    x"4F",x"06",x"00",x"21",x"6C",x"1F",x"09",x"4E", -- 0x0EE8
    x"2C",x"66",x"69",x"7E",x"0F",x"0F",x"D6",x"10", -- 0x0EF0
    x"4F",x"2C",x"2C",x"46",x"7A",x"93",x"D8",x"91", -- 0x0EF8
    x"38",x"02",x"10",x"F9",x"81",x"47",x"DD",x"6E", -- 0x0F00
    x"0B",x"26",x"80",x"7E",x"DD",x"77",x"02",x"90", -- 0x0F08
    x"DD",x"77",x"01",x"81",x"DD",x"77",x"00",x"CD", -- 0x0F10
    x"11",x"0B",x"0F",x"38",x"0A",x"DD",x"36",x"05", -- 0x0F18
    x"80",x"DD",x"36",x"03",x"F0",x"18",x"08",x"DD", -- 0x0F20
    x"36",x"05",x"00",x"DD",x"36",x"03",x"00",x"DD", -- 0x0F28
    x"36",x"06",x"01",x"DD",x"36",x"09",x"08",x"C9", -- 0x0F30
    x"DD",x"7E",x"06",x"B7",x"C8",x"DD",x"7E",x"04", -- 0x0F38
    x"21",x"47",x"80",x"BE",x"C0",x"DD",x"7E",x"05", -- 0x0F40
    x"B7",x"FD",x"7E",x"00",x"21",x"44",x"80",x"20", -- 0x0F48
    x"04",x"C6",x"14",x"18",x"02",x"D6",x"04",x"96", -- 0x0F50
    x"D8",x"FE",x"10",x"D0",x"3E",x"01",x"32",x"04", -- 0x0F58
    x"80",x"DD",x"36",x"06",x"02",x"C9",x"2C",x"2E", -- 0x0F60
    x"30",x"2E",x"27",x"38",x"70",x"82",x"73",x"82", -- 0x0F68
    x"76",x"82",x"79",x"82",x"7C",x"82",x"50",x"0C", -- 0x0F70
    x"30",x"10",x"70",x"14",x"40",x"18",x"40",x"1C", -- 0x0F78
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F80
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F88
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F90
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F98
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
