library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pace_pkg.all;
use work.kbd_pkg.all;

entity Game is
  port
  (
    -- clocking and reset
    clk							: in std_logic_vector(0 to 3);                       
    reset           : in std_logic;                       
    test_button     : in std_logic;                       

    -- inputs
    ps2clk          : inout std_logic;                       
    ps2data         : inout std_logic;                       
    dip             : in std_logic_vector(7 downto 0);    
		jamma						: in JAMMAInputsType;
		
    -- micro buses
    upaddr          : out std_logic_vector(15 downto 0);   
    updatao         : out std_logic_vector(7 downto 0);    

    -- SRAM
		sram_i					: in from_SRAM_t;
		sram_o					: out to_SRAM_t;

    gfxextra_data   : out std_logic_vector(7 downto 0);
		palette_data		: out ByteArrayType(15 downto 0);

    -- graphics (bitmap)
    bitmap_addr			: in std_logic_vector(15 downto 0);   
    bitmap_data			: out std_logic_vector(7 downto 0);    

    -- graphics (tilemap)
    tileaddr        : in std_logic_vector(15 downto 0);   
    tiledatao       : out std_logic_vector(7 downto 0);    
    tilemapaddr     : in std_logic_vector(15 downto 0);   
    tilemapdatao    : out std_logic_vector(15 downto 0);    
    attr_addr       : in std_logic_vector(9 downto 0);    
    attr_dout       : out std_logic_vector(15 downto 0);   

    -- graphics (sprite)
    sprite_reg_addr : out std_logic_vector(7 downto 0);    
    sprite_wr       : out std_logic;                       
    spriteaddr      : in std_logic_vector(15 downto 0);   
    spritedata      : out std_logic_vector(31 downto 0);
		spr0_hit				: in std_logic;

    -- graphics (control)
    vblank          : in std_logic;    
		xcentre					: out std_logic_vector(9 downto 0);
		ycentre					: out std_logic_vector(9 downto 0);

    -- OSD
    to_osd          : out to_OSD_t;
    from_osd        : in from_OSD_t;

    -- sound
    snd_rd          : out std_logic;                       
    snd_wr          : out std_logic;
    sndif_datai     : in std_logic_vector(7 downto 0);    

    -- spi interface
    spi_clk         : out std_logic;                       
    spi_din         : in std_logic;                       
    spi_dout        : out std_logic;                       
    spi_ena         : out std_logic;                       
    spi_mode        : out std_logic;                       
    spi_sel         : out std_logic;                       

    -- serial
    ser_rx          : in std_logic;                       
    ser_tx          : out std_logic;                       

    -- on-board leds
    leds            : out std_logic_vector(7 downto 0)    
  );
end Game;

architecture SYN of Game is

	alias clk_30M					: std_logic is clk(0);
	alias clk_40M					: std_logic is clk(1);
	
	signal reset_n				: std_logic;
	
  -- uP signals  
  signal clk_1M5_en			: std_logic;
  signal up_addr        : std_logic_vector(23 downto 0);
	alias addr_bus				: std_logic_vector(13 downto 0) is up_addr(13 downto 0);
  signal up_datai       : std_logic_vector(7 downto 0);
  signal up_datao       : std_logic_vector(7 downto 0);
  signal up_rw_n				: std_logic;
  signal up_irq_n				: std_logic;
	                        
  -- ROM signals        
	signal rom_cs					: std_logic;
  signal rom_data      	: std_logic_vector(7 downto 0);
                        
  -- keyboard signals
	                        
  -- VRAM signals       
	signal vram_cs				: std_logic;
	signal vram_wr				: std_logic;
	signal vram_addr			: std_logic_vector(9 downto 0);
  signal vram_datao     : std_logic_vector(7 downto 0);
                        
  -- RAM signals        
  signal wram_cs        : std_logic;
	signal wram_wr				: std_logic;
  alias wram_datao     	: std_logic_vector(7 downto 0) is sram_i.d(7 downto 0);

  -- RAM signals        
  signal cram_cs        : std_logic;
  signal cram_wr        : std_logic;
	signal cram0_wr				: std_logic;
	signal cram1_wr				: std_logic;
	signal cram0_datao		: std_logic_vector(7 downto 0);
	signal cram1_datao		: std_logic_vector(7 downto 0);
	
  -- other signals      
  signal dip_cs 				: std_logic;
  signal in0_cs 				: std_logic;
  signal in1_cs 				: std_logic;
  signal in2_cs 				: std_logic;
  signal in3_cs 				: std_logic;
	signal pokey_cs 			: std_logic;
  signal intack_wr			: std_logic;
	signal inputs					: in8(0 to 2);
	signal vblank_n				: std_logic;			-- should be vsync, but we don't have that
	signal vblank_fake		: std_logic;			-- generated by intgen, not video controller
	
	signal newtileAddr		: std_logic_vector(11 downto 0);
	
begin

	reset_n <= not reset;
	vblank_n <= not vblank;
	
	xcentre <= (others => '0');
	ycentre <= (others => '0');
	
  -- centipede A15 & A14 aren't connected on the PCB
  -- chip select logic

	-- WRAM $0000-$03FF
	-- SPRITE_RAM $07C0-$07FF (use SRAM atm)
	-- atari_vg_earom $1700-$173F
	wram_cs <= 	'1' when STD_MATCH(addr_bus, "0000----------") else 
							'1' when STD_MATCH(addr_bus, "00011111------") else
							'1' when STD_MATCH(addr_bus, "01011100------") else
							'0';
	-- VRAM $0400-$07BF
	vram_cs <= 	'1' when addr_bus(13 downto 10) = "0001" and addr_bus(9 downto 6) /= "1111" else '0';
	-- DIP0 $0800
  dip_cs <= 	'1' when STD_MATCH(addr_bus, "00100000000000") else '0';
	-- IN0 $0C00 (analog?)
  in0_cs <= 	'1' when STD_MATCH(addr_bus, "00110000000000") else '0';
	-- IN1 $0C01 (digital)
  in1_cs <= 	'1' when STD_MATCH(addr_bus, "00110000000001") else '0';
	-- IN2 $0C02 (analog?)
  in2_cs <= 	'1' when STD_MATCH(addr_bus, "00110000000010") else '0';
	-- IN3 $0C03 (digital)
  in3_cs <= 	'1' when STD_MATCH(addr_bus, "00110000000011") else '0';
	-- POKEY $1000-$100F
	pokey_cs <=	'1' when STD_MATCH(addr_bus, "0100000000----") else '0';
	-- ROM $2000-$3FFF
  rom_cs <= 	'1' when STD_MATCH(addr_bus, "1-------------") else '0';

	-- memory read mux
	uP_datai <= vram_datao when vram_cs = '1' else
							not dip when dip_cs = '1' else
							(inputs(0)(7) & vblank_fake & inputs(0)(5 downto 0)) when in0_cs = '1' else
							inputs(1) when in1_cs = '1' else
							inputs(2) when in2_cs = '1' else
							X"00" when in3_cs = '1' else
							sndif_datai when pokey_cs = '1' else
							rom_data when rom_cs = '1' else
							wram_datao;

  snd_rd <= up_rw_n and pokey_cs;

	-- wram $0000-$03FF
	-- sprite_wr $07C0-$07FF
	-- atari_vg_earom $1600-$163F
  -- atari_vg_earom_ctrl $1680
	-- * handled below
  -- vram_wr $0400-$07BF
	vram_wr <= not up_rw_n and vram_cs;
	-- sprite_wr $07C0-$07FF
  sprite_wr <= not up_rw_n when addr_bus(13 downto 6) = "00011111" else '0';
	-- POKEY $1000-$100F
  snd_wr <= not up_rw_n and pokey_cs;
	-- palette ram $1400-$140F
  cram_wr <= not up_rw_n when addr_bus(13 downto 4) = "0101000000" else '0';
	-- intack_wr $1800
  intack_wr <= not up_rw_n when addr_bus = "01100000000000" else '0';

  -- sprite register address
  -- sprite registers for sprite #0 @ $00,$10,$20,$30
  -- sprite registers for sprite #1 @ $01,$11,$21,$31
  sprite_reg_addr <= addr_bus(7 downto 6) & addr_bus(3 downto 0) & addr_bus(5 downto 4);

	-- mangle sprite address according to tile layout
	newTileAddr <= tileAddr(11 downto 5) & tileAddr(3 downto 1) & tileAddr(4) & tileAddr(0);

  -- SRAM signals (may or may not be used)
  sram_o.a <= std_logic_vector(resize(unsigned(addr_bus), sram_o.a'length));
  sram_o.d <= std_logic_vector(resize(unsigned(up_datao), sram_o.d'length));
	sram_o.be <= std_logic_vector(to_unsigned(1, sram_o.be'length));
  sram_o.cs <= '1';
  sram_o.oe <= wram_cs and up_rw_n;
  sram_o.we <= wram_cs and not up_rw_n;
	
	upaddr <= up_addr(upaddr'range);
	updatao <= up_datao;

  gfxextra_data <= (others => '0');
	GEN_PAL_DAT : for i in palette_data'range generate
		palette_data(i) <= (others => '0');
	end generate GEN_PAL_DAT;

  -- unused outputs
	bitmap_data <= (others => '0');
	spi_clk <= '0';
	spi_dout <= '0';
	spi_ena <= '0';
	spi_mode <= '0';
	spi_sel <= '0';
	ser_tx <= 'X';
	leds <= inputs(0);
	
  --
  -- COMPONENT INSTANTIATION
  --

	-- generate CPU clock enable (1M5Hz from 30MHz)
	clk_en_inst : entity work.clk_div
		generic map
		(
			DIVISOR		=> 20
		)
		port map
		(
			clk				=> clk_30M,
			reset			=> reset,
			clk_en		=> clk_1M5_en
		);

	up_inst : entity work.T65
		port map
		(
			Mode    		=> "00",	-- 6502
			Res_n   		=> reset_n,
			Enable  		=> clk_1M5_en,
			Clk     		=> clk_30M,
			Rdy     		=> '1',
			Abort_n 		=> '1',
			IRQ_n   		=> up_irq_n,
			NMI_n   		=> '1',
			SO_n    		=> '1',
			R_W_n   		=> up_rw_n,
			Sync    		=> open,
			EF      		=> open,
			MF      		=> open,
			XF      		=> open,
			ML_n    		=> open,
			VP_n    		=> open,
			VDA     		=> open,
			VPA     		=> open,
			A       		=> up_addr,
			DI      		=> up_datai,
			DO      		=> up_datao
		);

	rom_inst : entity work.sprom
		generic map
		(
			init_file		=> "../../../../src/platform/centiped/roms/rom0.hex",
			numwords_a	=> 8192,
			widthad_a		=> 13
		)
		port map
		(
			clock			=> clk_30M,
			address		=> addr_bus(12 downto 0),
			q					=> rom_data
		);
	
	vram_inst : entity work.dpram
		-- wren_a *MUST* be GND for CYCLONEII_SAFE_WRITE=VERIFIED_SAFE
		generic map
		(
			init_file		=> "../../../../src/platform/centiped/roms/vram.hex",
			numwords_a	=> 1024,
			widthad_a		=> 10
		)
		port map
		(
			clock_b			=> clk_30M,
			address_b		=> addr_bus(9 downto 0),
			wren_b			=> vram_wr,
			data_b			=> up_datao,
			q_b					=> vram_datao,

			clock_a			=> clk_40M,
			address_a		=> vram_addr,
			wren_a			=> '0',
			data_a			=> (others => 'X'),
			q_a					=> tileMapDatao(7 downto 0)
		);
	tilemapdatao(15 downto 8) <= (others => '0');
	
	vrammapper_inst : entity work.vramMapper
		port map
		(
	    clk     => clk_40M,

	    inAddr  => tileMapAddr(12 downto 0),
	    outAddr => vram_addr
		);

	cram0_wr <= cram_wr and not addr_bus(0);
	
	-- wren_a *MUST* be GND for CYCLONEII_SAFE_WRITE=VERIFIED_SAFE
	cram_inst_0 : entity work.dpram
		generic map
		(
			numwords_a			=> 128,
			widthad_a				=> 7
		)
		port map
		(
			clock_b					=> clk_30M,
			address_b				=> addr_bus(7 downto 1),
			wren_b					=> cram0_wr,
			data_b					=> up_datao,
			q_b							=> cram0_datao,
			
			clock_a					=> clk_40M,
			address_a				=> attr_addr(7 downto 1),
			wren_a					=> '0',
			data_a					=> (others => 'X'),
			q_a							=> attr_dout(7 downto 0)
		);

	cram1_wr <= cram_wr and addr_bus(0);

	-- wren_a *MUST* be GND for CYCLONEII_SAFE_WRITE=VERIFIED_SAFE
	cram_inst_1 : entity work.dpram
		generic map
		(
			numwords_a			=> 128,
			widthad_a				=> 7
		)
		port map
		(
			clock_b					=> clk_30M,
			address_b				=> addr_bus(7 downto 1),
			wren_b					=> cram1_wr,
			data_b					=> up_datao,
			q_b							=> cram1_datao,
			
			clock_a					=> clk_40M,
			address_a				=> attr_addr(7 downto 1),
			wren_a					=> '0',
			data_a					=> (others => 'X'),
			q_a							=> attr_dout(15 downto 8)
		);

	inputs_inst : entity work.Inputs
		generic map
		(
			NUM_INPUTS	=> 3
		)
	  port map
	  (
	    clk     		=> clk_30M,
	    reset   		=> reset,
	    ps2clk  		=> ps2clk,
	    ps2data 		=> ps2data,
			jamma				=> jamma,

	    dips				=> dip,
	    inputs			=> inputs
	  );

	intgen_inst : entity work.intGen
		port map
		(
	    clk       	=> clk_30M,
	    reset     	=> reset,

	    -- inputs
	    vsync_n   	=> vblank_n,
	    intack    	=> intack_wr,

	    -- outputs
	    vblank    	=> vblank_fake,
	    irq_n     	=> up_irq_n
		);

	gfxrom_inst : entity work.dprom_2r
		generic map
		(
			init_file		=> "../../../../src/platform/centiped/roms/gfxrom.hex",
			numwords_a	=> 4096,
			widthad_a		=> 12,
			numwords_b	=> 1024,
			widthad_b		=> 10,
			width_b			=> 32
		)
		port map
		(
			clock										=> clk_40M,
			address_a								=> newtileaddr(11 downto 0),
			q_a											=> tileDatao,
			
			address_b								=> spriteaddr(9 downto 0),
			q_b(31 downto 24)				=> spriteData(7 downto 0),
			q_b(23 downto 16)				=> spriteData(15 downto 8),
			q_b(15 downto 8)				=> spriteData(23 downto 16),
			q_b(7 downto 0)					=> spriteData(31 downto 24)
		);

end SYN;
