-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VIC20_BASIC_ROM is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of VIC20_BASIC_ROM is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"78",x"E3",x"67",x"E4",x"43",x"42",x"4D",x"42", -- 0x0000
    x"41",x"53",x"49",x"43",x"30",x"C8",x"41",x"C7", -- 0x0008
    x"1D",x"CD",x"F7",x"C8",x"A4",x"CB",x"BE",x"CB", -- 0x0010
    x"80",x"D0",x"05",x"CC",x"A4",x"C9",x"9F",x"C8", -- 0x0018
    x"70",x"C8",x"27",x"C9",x"1C",x"C8",x"82",x"C8", -- 0x0020
    x"D1",x"C8",x"3A",x"C9",x"2E",x"C8",x"4A",x"C9", -- 0x0028
    x"2C",x"D8",x"64",x"E1",x"52",x"E1",x"61",x"E1", -- 0x0030
    x"B2",x"D3",x"23",x"D8",x"7F",x"CA",x"9F",x"CA", -- 0x0038
    x"56",x"C8",x"9B",x"C6",x"5D",x"C6",x"85",x"CA", -- 0x0040
    x"26",x"E1",x"BA",x"E1",x"C3",x"E1",x"7A",x"CB", -- 0x0048
    x"41",x"C6",x"39",x"DC",x"CC",x"DC",x"58",x"DC", -- 0x0050
    x"00",x"00",x"7D",x"D3",x"9E",x"D3",x"71",x"DF", -- 0x0058
    x"94",x"E0",x"EA",x"D9",x"ED",x"DF",x"61",x"E2", -- 0x0060
    x"68",x"E2",x"B1",x"E2",x"0B",x"E3",x"0D",x"D8", -- 0x0068
    x"7C",x"D7",x"65",x"D4",x"AD",x"D7",x"8B",x"D7", -- 0x0070
    x"EC",x"D6",x"00",x"D7",x"2C",x"D7",x"37",x"D7", -- 0x0078
    x"79",x"69",x"D8",x"79",x"52",x"D8",x"7B",x"2A", -- 0x0080
    x"DA",x"7B",x"11",x"DB",x"7F",x"7A",x"DF",x"50", -- 0x0088
    x"E8",x"CF",x"46",x"E5",x"CF",x"7D",x"B3",x"DF", -- 0x0090
    x"5A",x"D3",x"CE",x"64",x"15",x"D0",x"45",x"4E", -- 0x0098
    x"C4",x"46",x"4F",x"D2",x"4E",x"45",x"58",x"D4", -- 0x00A0
    x"44",x"41",x"54",x"C1",x"49",x"4E",x"50",x"55", -- 0x00A8
    x"54",x"A3",x"49",x"4E",x"50",x"55",x"D4",x"44", -- 0x00B0
    x"49",x"CD",x"52",x"45",x"41",x"C4",x"4C",x"45", -- 0x00B8
    x"D4",x"47",x"4F",x"54",x"CF",x"52",x"55",x"CE", -- 0x00C0
    x"49",x"C6",x"52",x"45",x"53",x"54",x"4F",x"52", -- 0x00C8
    x"C5",x"47",x"4F",x"53",x"55",x"C2",x"52",x"45", -- 0x00D0
    x"54",x"55",x"52",x"CE",x"52",x"45",x"CD",x"53", -- 0x00D8
    x"54",x"4F",x"D0",x"4F",x"CE",x"57",x"41",x"49", -- 0x00E0
    x"D4",x"4C",x"4F",x"41",x"C4",x"53",x"41",x"56", -- 0x00E8
    x"C5",x"56",x"45",x"52",x"49",x"46",x"D9",x"44", -- 0x00F0
    x"45",x"C6",x"50",x"4F",x"4B",x"C5",x"50",x"52", -- 0x00F8
    x"49",x"4E",x"54",x"A3",x"50",x"52",x"49",x"4E", -- 0x0100
    x"D4",x"43",x"4F",x"4E",x"D4",x"4C",x"49",x"53", -- 0x0108
    x"D4",x"43",x"4C",x"D2",x"43",x"4D",x"C4",x"53", -- 0x0110
    x"59",x"D3",x"4F",x"50",x"45",x"CE",x"43",x"4C", -- 0x0118
    x"4F",x"53",x"C5",x"47",x"45",x"D4",x"4E",x"45", -- 0x0120
    x"D7",x"54",x"41",x"42",x"A8",x"54",x"CF",x"46", -- 0x0128
    x"CE",x"53",x"50",x"43",x"A8",x"54",x"48",x"45", -- 0x0130
    x"CE",x"4E",x"4F",x"D4",x"53",x"54",x"45",x"D0", -- 0x0138
    x"AB",x"AD",x"AA",x"AF",x"DE",x"41",x"4E",x"C4", -- 0x0140
    x"4F",x"D2",x"BE",x"BD",x"BC",x"53",x"47",x"CE", -- 0x0148
    x"49",x"4E",x"D4",x"41",x"42",x"D3",x"55",x"53", -- 0x0150
    x"D2",x"46",x"52",x"C5",x"50",x"4F",x"D3",x"53", -- 0x0158
    x"51",x"D2",x"52",x"4E",x"C4",x"4C",x"4F",x"C7", -- 0x0160
    x"45",x"58",x"D0",x"43",x"4F",x"D3",x"53",x"49", -- 0x0168
    x"CE",x"54",x"41",x"CE",x"41",x"54",x"CE",x"50", -- 0x0170
    x"45",x"45",x"CB",x"4C",x"45",x"CE",x"53",x"54", -- 0x0178
    x"52",x"A4",x"56",x"41",x"CC",x"41",x"53",x"C3", -- 0x0180
    x"43",x"48",x"52",x"A4",x"4C",x"45",x"46",x"54", -- 0x0188
    x"A4",x"52",x"49",x"47",x"48",x"54",x"A4",x"4D", -- 0x0190
    x"49",x"44",x"A4",x"47",x"CF",x"00",x"54",x"4F", -- 0x0198
    x"4F",x"20",x"4D",x"41",x"4E",x"59",x"20",x"46", -- 0x01A0
    x"49",x"4C",x"45",x"D3",x"46",x"49",x"4C",x"45", -- 0x01A8
    x"20",x"4F",x"50",x"45",x"CE",x"46",x"49",x"4C", -- 0x01B0
    x"45",x"20",x"4E",x"4F",x"54",x"20",x"4F",x"50", -- 0x01B8
    x"45",x"CE",x"46",x"49",x"4C",x"45",x"20",x"4E", -- 0x01C0
    x"4F",x"54",x"20",x"46",x"4F",x"55",x"4E",x"C4", -- 0x01C8
    x"44",x"45",x"56",x"49",x"43",x"45",x"20",x"4E", -- 0x01D0
    x"4F",x"54",x"20",x"50",x"52",x"45",x"53",x"45", -- 0x01D8
    x"4E",x"D4",x"4E",x"4F",x"54",x"20",x"49",x"4E", -- 0x01E0
    x"50",x"55",x"54",x"20",x"46",x"49",x"4C",x"C5", -- 0x01E8
    x"4E",x"4F",x"54",x"20",x"4F",x"55",x"54",x"50", -- 0x01F0
    x"55",x"54",x"20",x"46",x"49",x"4C",x"C5",x"4D", -- 0x01F8
    x"49",x"53",x"53",x"49",x"4E",x"47",x"20",x"46", -- 0x0200
    x"49",x"4C",x"45",x"20",x"4E",x"41",x"4D",x"C5", -- 0x0208
    x"49",x"4C",x"4C",x"45",x"47",x"41",x"4C",x"20", -- 0x0210
    x"44",x"45",x"56",x"49",x"43",x"45",x"20",x"4E", -- 0x0218
    x"55",x"4D",x"42",x"45",x"D2",x"4E",x"45",x"58", -- 0x0220
    x"54",x"20",x"57",x"49",x"54",x"48",x"4F",x"55", -- 0x0228
    x"54",x"20",x"46",x"4F",x"D2",x"53",x"59",x"4E", -- 0x0230
    x"54",x"41",x"D8",x"52",x"45",x"54",x"55",x"52", -- 0x0238
    x"4E",x"20",x"57",x"49",x"54",x"48",x"4F",x"55", -- 0x0240
    x"54",x"20",x"47",x"4F",x"53",x"55",x"C2",x"4F", -- 0x0248
    x"55",x"54",x"20",x"4F",x"46",x"20",x"44",x"41", -- 0x0250
    x"54",x"C1",x"49",x"4C",x"4C",x"45",x"47",x"41", -- 0x0258
    x"4C",x"20",x"51",x"55",x"41",x"4E",x"54",x"49", -- 0x0260
    x"54",x"D9",x"4F",x"56",x"45",x"52",x"46",x"4C", -- 0x0268
    x"4F",x"D7",x"4F",x"55",x"54",x"20",x"4F",x"46", -- 0x0270
    x"20",x"4D",x"45",x"4D",x"4F",x"52",x"D9",x"55", -- 0x0278
    x"4E",x"44",x"45",x"46",x"27",x"44",x"20",x"53", -- 0x0280
    x"54",x"41",x"54",x"45",x"4D",x"45",x"4E",x"D4", -- 0x0288
    x"42",x"41",x"44",x"20",x"53",x"55",x"42",x"53", -- 0x0290
    x"43",x"52",x"49",x"50",x"D4",x"52",x"45",x"44", -- 0x0298
    x"49",x"4D",x"27",x"44",x"20",x"41",x"52",x"52", -- 0x02A0
    x"41",x"D9",x"44",x"49",x"56",x"49",x"53",x"49", -- 0x02A8
    x"4F",x"4E",x"20",x"42",x"59",x"20",x"5A",x"45", -- 0x02B0
    x"52",x"CF",x"49",x"4C",x"4C",x"45",x"47",x"41", -- 0x02B8
    x"4C",x"20",x"44",x"49",x"52",x"45",x"43",x"D4", -- 0x02C0
    x"54",x"59",x"50",x"45",x"20",x"4D",x"49",x"53", -- 0x02C8
    x"4D",x"41",x"54",x"43",x"C8",x"53",x"54",x"52", -- 0x02D0
    x"49",x"4E",x"47",x"20",x"54",x"4F",x"4F",x"20", -- 0x02D8
    x"4C",x"4F",x"4E",x"C7",x"46",x"49",x"4C",x"45", -- 0x02E0
    x"20",x"44",x"41",x"54",x"C1",x"46",x"4F",x"52", -- 0x02E8
    x"4D",x"55",x"4C",x"41",x"20",x"54",x"4F",x"4F", -- 0x02F0
    x"20",x"43",x"4F",x"4D",x"50",x"4C",x"45",x"D8", -- 0x02F8
    x"43",x"41",x"4E",x"27",x"54",x"20",x"43",x"4F", -- 0x0300
    x"4E",x"54",x"49",x"4E",x"55",x"C5",x"55",x"4E", -- 0x0308
    x"44",x"45",x"46",x"27",x"44",x"20",x"46",x"55", -- 0x0310
    x"4E",x"43",x"54",x"49",x"4F",x"CE",x"56",x"45", -- 0x0318
    x"52",x"49",x"46",x"D9",x"4C",x"4F",x"41",x"C4", -- 0x0320
    x"9E",x"C1",x"AC",x"C1",x"B5",x"C1",x"C2",x"C1", -- 0x0328
    x"D0",x"C1",x"E2",x"C1",x"F0",x"C1",x"FF",x"C1", -- 0x0330
    x"10",x"C2",x"25",x"C2",x"35",x"C2",x"3B",x"C2", -- 0x0338
    x"4F",x"C2",x"5A",x"C2",x"6A",x"C2",x"72",x"C2", -- 0x0340
    x"7F",x"C2",x"90",x"C2",x"9D",x"C2",x"AA",x"C2", -- 0x0348
    x"BA",x"C2",x"C8",x"C2",x"D5",x"C2",x"E4",x"C2", -- 0x0350
    x"ED",x"C2",x"00",x"C3",x"0E",x"C3",x"1E",x"C3", -- 0x0358
    x"24",x"C3",x"83",x"C3",x"0D",x"4F",x"4B",x"0D", -- 0x0360
    x"00",x"0D",x"20",x"45",x"52",x"52",x"4F",x"52", -- 0x0368
    x"00",x"20",x"49",x"4E",x"20",x"00",x"0D",x"0A", -- 0x0370
    x"52",x"45",x"41",x"44",x"59",x"2E",x"0D",x"0A", -- 0x0378
    x"00",x"0D",x"0A",x"42",x"52",x"45",x"41",x"4B", -- 0x0380
    x"00",x"A0",x"BA",x"E8",x"E8",x"E8",x"E8",x"BD", -- 0x0388
    x"01",x"01",x"C9",x"81",x"D0",x"21",x"A5",x"4A", -- 0x0390
    x"D0",x"0A",x"BD",x"02",x"01",x"85",x"49",x"BD", -- 0x0398
    x"03",x"01",x"85",x"4A",x"DD",x"03",x"01",x"D0", -- 0x03A0
    x"07",x"A5",x"49",x"DD",x"02",x"01",x"F0",x"07", -- 0x03A8
    x"8A",x"18",x"69",x"12",x"AA",x"D0",x"D8",x"60", -- 0x03B0
    x"20",x"08",x"C4",x"85",x"31",x"84",x"32",x"38", -- 0x03B8
    x"A5",x"5A",x"E5",x"5F",x"85",x"22",x"A8",x"A5", -- 0x03C0
    x"5B",x"E5",x"60",x"AA",x"E8",x"98",x"F0",x"23", -- 0x03C8
    x"A5",x"5A",x"38",x"E5",x"22",x"85",x"5A",x"B0", -- 0x03D0
    x"03",x"C6",x"5B",x"38",x"A5",x"58",x"E5",x"22", -- 0x03D8
    x"85",x"58",x"B0",x"08",x"C6",x"59",x"90",x"04", -- 0x03E0
    x"B1",x"5A",x"91",x"58",x"88",x"D0",x"F9",x"B1", -- 0x03E8
    x"5A",x"91",x"58",x"C6",x"5B",x"C6",x"59",x"CA", -- 0x03F0
    x"D0",x"F2",x"60",x"0A",x"69",x"3E",x"B0",x"35", -- 0x03F8
    x"85",x"22",x"BA",x"E4",x"22",x"90",x"2E",x"60", -- 0x0400
    x"C4",x"34",x"90",x"28",x"D0",x"04",x"C5",x"33", -- 0x0408
    x"90",x"22",x"48",x"A2",x"09",x"98",x"48",x"B5", -- 0x0410
    x"57",x"CA",x"10",x"FA",x"20",x"26",x"D5",x"A2", -- 0x0418
    x"F7",x"68",x"95",x"61",x"E8",x"30",x"FA",x"68", -- 0x0420
    x"A8",x"68",x"C4",x"34",x"90",x"06",x"D0",x"05", -- 0x0428
    x"C5",x"33",x"B0",x"01",x"60",x"A2",x"10",x"6C", -- 0x0430
    x"00",x"03",x"8A",x"0A",x"AA",x"BD",x"26",x"C3", -- 0x0438
    x"85",x"22",x"BD",x"27",x"C3",x"85",x"23",x"20", -- 0x0440
    x"CC",x"FF",x"A9",x"00",x"85",x"13",x"20",x"D7", -- 0x0448
    x"CA",x"20",x"45",x"CB",x"A0",x"00",x"B1",x"22", -- 0x0450
    x"48",x"29",x"7F",x"20",x"47",x"CB",x"C8",x"68", -- 0x0458
    x"10",x"F4",x"20",x"7A",x"C6",x"A9",x"69",x"A0", -- 0x0460
    x"C3",x"20",x"1E",x"CB",x"A4",x"3A",x"C8",x"F0", -- 0x0468
    x"03",x"20",x"C2",x"DD",x"A9",x"76",x"A0",x"C3", -- 0x0470
    x"20",x"1E",x"CB",x"A9",x"80",x"20",x"90",x"FF", -- 0x0478
    x"6C",x"02",x"03",x"20",x"60",x"C5",x"86",x"7A", -- 0x0480
    x"84",x"7B",x"20",x"73",x"00",x"AA",x"F0",x"F0", -- 0x0488
    x"A2",x"FF",x"86",x"3A",x"90",x"06",x"20",x"79", -- 0x0490
    x"C5",x"4C",x"E1",x"C7",x"20",x"6B",x"C9",x"20", -- 0x0498
    x"79",x"C5",x"84",x"0B",x"20",x"13",x"C6",x"90", -- 0x04A0
    x"44",x"A0",x"01",x"B1",x"5F",x"85",x"23",x"A5", -- 0x04A8
    x"2D",x"85",x"22",x"A5",x"60",x"85",x"25",x"A5", -- 0x04B0
    x"5F",x"88",x"F1",x"5F",x"18",x"65",x"2D",x"85", -- 0x04B8
    x"2D",x"85",x"24",x"A5",x"2E",x"69",x"FF",x"85", -- 0x04C0
    x"2E",x"E5",x"60",x"AA",x"38",x"A5",x"5F",x"E5", -- 0x04C8
    x"2D",x"A8",x"B0",x"03",x"E8",x"C6",x"25",x"18", -- 0x04D0
    x"65",x"22",x"90",x"03",x"C6",x"23",x"18",x"B1", -- 0x04D8
    x"22",x"91",x"24",x"C8",x"D0",x"F9",x"E6",x"23", -- 0x04E0
    x"E6",x"25",x"CA",x"D0",x"F2",x"20",x"59",x"C6", -- 0x04E8
    x"20",x"33",x"C5",x"AD",x"00",x"02",x"F0",x"88", -- 0x04F0
    x"18",x"A5",x"2D",x"85",x"5A",x"65",x"0B",x"85", -- 0x04F8
    x"58",x"A4",x"2E",x"84",x"5B",x"90",x"01",x"C8", -- 0x0500
    x"84",x"59",x"20",x"B8",x"C3",x"A5",x"14",x"A4", -- 0x0508
    x"15",x"8D",x"FE",x"01",x"8C",x"FF",x"01",x"A5", -- 0x0510
    x"31",x"A4",x"32",x"85",x"2D",x"84",x"2E",x"A4", -- 0x0518
    x"0B",x"88",x"B9",x"FC",x"01",x"91",x"5F",x"88", -- 0x0520
    x"10",x"F8",x"20",x"59",x"C6",x"20",x"33",x"C5", -- 0x0528
    x"4C",x"80",x"C4",x"A5",x"2B",x"A4",x"2C",x"85", -- 0x0530
    x"22",x"84",x"23",x"18",x"A0",x"01",x"B1",x"22", -- 0x0538
    x"F0",x"1D",x"A0",x"04",x"C8",x"B1",x"22",x"D0", -- 0x0540
    x"FB",x"C8",x"98",x"65",x"22",x"AA",x"A0",x"00", -- 0x0548
    x"91",x"22",x"A5",x"23",x"69",x"00",x"C8",x"91", -- 0x0550
    x"22",x"86",x"22",x"85",x"23",x"90",x"DD",x"60", -- 0x0558
    x"A2",x"00",x"20",x"0F",x"E1",x"C9",x"0D",x"F0", -- 0x0560
    x"0D",x"9D",x"00",x"02",x"E8",x"E0",x"59",x"90", -- 0x0568
    x"F1",x"A2",x"17",x"4C",x"37",x"C4",x"4C",x"CA", -- 0x0570
    x"CA",x"6C",x"04",x"03",x"A6",x"7A",x"A0",x"04", -- 0x0578
    x"84",x"0F",x"BD",x"00",x"02",x"10",x"07",x"C9", -- 0x0580
    x"FF",x"F0",x"3E",x"E8",x"D0",x"F4",x"C9",x"20", -- 0x0588
    x"F0",x"37",x"85",x"08",x"C9",x"22",x"F0",x"56", -- 0x0590
    x"24",x"0F",x"70",x"2D",x"C9",x"3F",x"D0",x"04", -- 0x0598
    x"A9",x"99",x"D0",x"25",x"C9",x"30",x"90",x"04", -- 0x05A0
    x"C9",x"3C",x"90",x"1D",x"84",x"71",x"A0",x"00", -- 0x05A8
    x"84",x"0B",x"88",x"86",x"7A",x"CA",x"C8",x"E8", -- 0x05B0
    x"BD",x"00",x"02",x"38",x"F9",x"9E",x"C0",x"F0", -- 0x05B8
    x"F5",x"C9",x"80",x"D0",x"30",x"05",x"0B",x"A4", -- 0x05C0
    x"71",x"E8",x"C8",x"99",x"FB",x"01",x"B9",x"FB", -- 0x05C8
    x"01",x"F0",x"36",x"38",x"E9",x"3A",x"F0",x"04", -- 0x05D0
    x"C9",x"49",x"D0",x"02",x"85",x"0F",x"38",x"E9", -- 0x05D8
    x"55",x"D0",x"9F",x"85",x"08",x"BD",x"00",x"02", -- 0x05E0
    x"F0",x"DF",x"C5",x"08",x"F0",x"DB",x"C8",x"99", -- 0x05E8
    x"FB",x"01",x"E8",x"D0",x"F0",x"A6",x"7A",x"E6", -- 0x05F0
    x"0B",x"C8",x"B9",x"9D",x"C0",x"10",x"FA",x"B9", -- 0x05F8
    x"9E",x"C0",x"D0",x"B4",x"BD",x"00",x"02",x"10", -- 0x0600
    x"BE",x"99",x"FD",x"01",x"C6",x"7B",x"A9",x"FF", -- 0x0608
    x"85",x"7A",x"60",x"A5",x"2B",x"A6",x"2C",x"A0", -- 0x0610
    x"01",x"85",x"5F",x"86",x"60",x"B1",x"5F",x"F0", -- 0x0618
    x"1F",x"C8",x"C8",x"A5",x"15",x"D1",x"5F",x"90", -- 0x0620
    x"18",x"F0",x"03",x"88",x"D0",x"09",x"A5",x"14", -- 0x0628
    x"88",x"D1",x"5F",x"90",x"0C",x"F0",x"0A",x"88", -- 0x0630
    x"B1",x"5F",x"AA",x"88",x"B1",x"5F",x"B0",x"D7", -- 0x0638
    x"18",x"60",x"D0",x"FD",x"A9",x"00",x"A8",x"91", -- 0x0640
    x"2B",x"C8",x"91",x"2B",x"A5",x"2B",x"18",x"69", -- 0x0648
    x"02",x"85",x"2D",x"A5",x"2C",x"69",x"00",x"85", -- 0x0650
    x"2E",x"20",x"8E",x"C6",x"A9",x"00",x"D0",x"2D", -- 0x0658
    x"20",x"E7",x"FF",x"A5",x"37",x"A4",x"38",x"85", -- 0x0660
    x"33",x"84",x"34",x"A5",x"2D",x"A4",x"2E",x"85", -- 0x0668
    x"2F",x"84",x"30",x"85",x"31",x"84",x"32",x"20", -- 0x0670
    x"1D",x"C8",x"A2",x"19",x"86",x"16",x"68",x"A8", -- 0x0678
    x"68",x"A2",x"FA",x"9A",x"48",x"98",x"48",x"A9", -- 0x0680
    x"00",x"85",x"3E",x"85",x"10",x"60",x"18",x"A5", -- 0x0688
    x"2B",x"69",x"FF",x"85",x"7A",x"A5",x"2C",x"69", -- 0x0690
    x"FF",x"85",x"7B",x"60",x"90",x"06",x"F0",x"04", -- 0x0698
    x"C9",x"AB",x"D0",x"E9",x"20",x"6B",x"C9",x"20", -- 0x06A0
    x"13",x"C6",x"20",x"79",x"00",x"F0",x"0C",x"C9", -- 0x06A8
    x"AB",x"D0",x"8E",x"20",x"73",x"00",x"20",x"6B", -- 0x06B0
    x"C9",x"D0",x"86",x"68",x"68",x"A5",x"14",x"05", -- 0x06B8
    x"15",x"D0",x"06",x"A9",x"FF",x"85",x"14",x"85", -- 0x06C0
    x"15",x"A0",x"01",x"84",x"0F",x"B1",x"5F",x"F0", -- 0x06C8
    x"43",x"20",x"2C",x"C8",x"20",x"D7",x"CA",x"C8", -- 0x06D0
    x"B1",x"5F",x"AA",x"C8",x"B1",x"5F",x"C5",x"15", -- 0x06D8
    x"D0",x"04",x"E4",x"14",x"F0",x"02",x"B0",x"2C", -- 0x06E0
    x"84",x"49",x"20",x"CD",x"DD",x"A9",x"20",x"A4", -- 0x06E8
    x"49",x"29",x"7F",x"20",x"47",x"CB",x"C9",x"22", -- 0x06F0
    x"D0",x"06",x"A5",x"0F",x"49",x"FF",x"85",x"0F", -- 0x06F8
    x"C8",x"F0",x"11",x"B1",x"5F",x"D0",x"10",x"A8", -- 0x0700
    x"B1",x"5F",x"AA",x"C8",x"B1",x"5F",x"86",x"5F", -- 0x0708
    x"85",x"60",x"D0",x"B5",x"4C",x"74",x"C4",x"6C", -- 0x0710
    x"06",x"03",x"10",x"D7",x"C9",x"FF",x"F0",x"D3", -- 0x0718
    x"24",x"0F",x"30",x"CF",x"38",x"E9",x"7F",x"AA", -- 0x0720
    x"84",x"49",x"A0",x"FF",x"CA",x"F0",x"08",x"C8", -- 0x0728
    x"B9",x"9E",x"C0",x"10",x"FA",x"30",x"F5",x"C8", -- 0x0730
    x"B9",x"9E",x"C0",x"30",x"B2",x"20",x"47",x"CB", -- 0x0738
    x"D0",x"F5",x"A9",x"80",x"85",x"10",x"20",x"A5", -- 0x0740
    x"C9",x"20",x"8A",x"C3",x"D0",x"05",x"8A",x"69", -- 0x0748
    x"0F",x"AA",x"9A",x"68",x"68",x"A9",x"09",x"20", -- 0x0750
    x"FB",x"C3",x"20",x"06",x"C9",x"18",x"98",x"65", -- 0x0758
    x"7A",x"48",x"A5",x"7B",x"69",x"00",x"48",x"A5", -- 0x0760
    x"3A",x"48",x"A5",x"39",x"48",x"A9",x"A4",x"20", -- 0x0768
    x"FF",x"CE",x"20",x"8D",x"CD",x"20",x"8A",x"CD", -- 0x0770
    x"A5",x"66",x"09",x"7F",x"25",x"62",x"85",x"62", -- 0x0778
    x"A9",x"8B",x"A0",x"C7",x"85",x"22",x"84",x"23", -- 0x0780
    x"4C",x"43",x"CE",x"A9",x"BC",x"A0",x"D9",x"20", -- 0x0788
    x"A2",x"DB",x"20",x"79",x"00",x"C9",x"A9",x"D0", -- 0x0790
    x"06",x"20",x"73",x"00",x"20",x"8A",x"CD",x"20", -- 0x0798
    x"2B",x"DC",x"20",x"38",x"CE",x"A5",x"4A",x"48", -- 0x07A0
    x"A5",x"49",x"48",x"A9",x"81",x"48",x"20",x"2C", -- 0x07A8
    x"C8",x"A5",x"7A",x"A4",x"7B",x"C0",x"02",x"EA", -- 0x07B0
    x"F0",x"04",x"85",x"3D",x"84",x"3E",x"A0",x"00", -- 0x07B8
    x"B1",x"7A",x"D0",x"43",x"A0",x"02",x"B1",x"7A", -- 0x07C0
    x"18",x"D0",x"03",x"4C",x"4B",x"C8",x"C8",x"B1", -- 0x07C8
    x"7A",x"85",x"39",x"C8",x"B1",x"7A",x"85",x"3A", -- 0x07D0
    x"98",x"65",x"7A",x"85",x"7A",x"90",x"02",x"E6", -- 0x07D8
    x"7B",x"6C",x"08",x"03",x"20",x"73",x"00",x"20", -- 0x07E0
    x"ED",x"C7",x"4C",x"AE",x"C7",x"F0",x"3C",x"E9", -- 0x07E8
    x"80",x"90",x"11",x"C9",x"23",x"B0",x"17",x"0A", -- 0x07F0
    x"A8",x"B9",x"0D",x"C0",x"48",x"B9",x"0C",x"C0", -- 0x07F8
    x"48",x"4C",x"73",x"00",x"4C",x"A5",x"C9",x"C9", -- 0x0800
    x"3A",x"F0",x"D6",x"4C",x"08",x"CF",x"C9",x"4B", -- 0x0808
    x"D0",x"F9",x"20",x"73",x"00",x"A9",x"A4",x"20", -- 0x0810
    x"FF",x"CE",x"4C",x"A0",x"C8",x"38",x"A5",x"2B", -- 0x0818
    x"E9",x"01",x"A4",x"2C",x"B0",x"01",x"88",x"85", -- 0x0820
    x"41",x"84",x"42",x"60",x"20",x"E1",x"FF",x"B0", -- 0x0828
    x"01",x"18",x"D0",x"3C",x"A5",x"7A",x"A4",x"7B", -- 0x0830
    x"A6",x"3A",x"E8",x"F0",x"0C",x"85",x"3D",x"84", -- 0x0838
    x"3E",x"A5",x"39",x"A4",x"3A",x"85",x"3B",x"84", -- 0x0840
    x"3C",x"68",x"68",x"A9",x"81",x"A0",x"C3",x"90", -- 0x0848
    x"03",x"4C",x"69",x"C4",x"4C",x"74",x"C4",x"D0", -- 0x0850
    x"17",x"A2",x"1A",x"A4",x"3E",x"D0",x"03",x"4C", -- 0x0858
    x"37",x"C4",x"A5",x"3D",x"85",x"7A",x"84",x"7B", -- 0x0860
    x"A5",x"3B",x"A4",x"3C",x"85",x"39",x"84",x"3A", -- 0x0868
    x"60",x"08",x"A9",x"00",x"20",x"90",x"FF",x"28", -- 0x0870
    x"D0",x"03",x"4C",x"59",x"C6",x"20",x"60",x"C6", -- 0x0878
    x"4C",x"97",x"C8",x"A9",x"03",x"20",x"FB",x"C3", -- 0x0880
    x"A5",x"7B",x"48",x"A5",x"7A",x"48",x"A5",x"3A", -- 0x0888
    x"48",x"A5",x"39",x"48",x"A9",x"8D",x"48",x"20", -- 0x0890
    x"79",x"00",x"20",x"A0",x"C8",x"4C",x"AE",x"C7", -- 0x0898
    x"20",x"6B",x"C9",x"20",x"09",x"C9",x"38",x"A5", -- 0x08A0
    x"39",x"E5",x"14",x"A5",x"3A",x"E5",x"15",x"B0", -- 0x08A8
    x"0B",x"98",x"38",x"65",x"7A",x"A6",x"7B",x"90", -- 0x08B0
    x"07",x"E8",x"B0",x"04",x"A5",x"2B",x"A6",x"2C", -- 0x08B8
    x"20",x"17",x"C6",x"90",x"1E",x"A5",x"5F",x"E9", -- 0x08C0
    x"01",x"85",x"7A",x"A5",x"60",x"E9",x"00",x"85", -- 0x08C8
    x"7B",x"60",x"D0",x"FD",x"A9",x"FF",x"85",x"4A", -- 0x08D0
    x"20",x"8A",x"C3",x"9A",x"C9",x"8D",x"F0",x"0B", -- 0x08D8
    x"A2",x"0C",x"2C",x"A2",x"11",x"4C",x"37",x"C4", -- 0x08E0
    x"4C",x"08",x"CF",x"68",x"68",x"85",x"39",x"68", -- 0x08E8
    x"85",x"3A",x"68",x"85",x"7A",x"68",x"85",x"7B", -- 0x08F0
    x"20",x"06",x"C9",x"98",x"18",x"65",x"7A",x"85", -- 0x08F8
    x"7A",x"90",x"02",x"E6",x"7B",x"60",x"A2",x"3A", -- 0x0900
    x"2C",x"A2",x"00",x"86",x"07",x"A0",x"00",x"84", -- 0x0908
    x"08",x"A5",x"08",x"A6",x"07",x"85",x"07",x"86", -- 0x0910
    x"08",x"B1",x"7A",x"F0",x"E8",x"C5",x"08",x"F0", -- 0x0918
    x"E4",x"C8",x"C9",x"22",x"D0",x"F3",x"F0",x"E9", -- 0x0920
    x"20",x"9E",x"CD",x"20",x"79",x"00",x"C9",x"89", -- 0x0928
    x"F0",x"05",x"A9",x"A7",x"20",x"FF",x"CE",x"A5", -- 0x0930
    x"61",x"D0",x"05",x"20",x"09",x"C9",x"F0",x"BB", -- 0x0938
    x"20",x"79",x"00",x"B0",x"03",x"4C",x"A0",x"C8", -- 0x0940
    x"4C",x"ED",x"C7",x"20",x"9E",x"D7",x"48",x"C9", -- 0x0948
    x"8D",x"F0",x"04",x"C9",x"89",x"D0",x"91",x"C6", -- 0x0950
    x"65",x"D0",x"04",x"68",x"4C",x"EF",x"C7",x"20", -- 0x0958
    x"73",x"00",x"20",x"6B",x"C9",x"C9",x"2C",x"F0", -- 0x0960
    x"EE",x"68",x"60",x"A2",x"00",x"86",x"14",x"86", -- 0x0968
    x"15",x"B0",x"F7",x"E9",x"2F",x"85",x"07",x"A5", -- 0x0970
    x"15",x"85",x"22",x"C9",x"19",x"B0",x"D4",x"A5", -- 0x0978
    x"14",x"0A",x"26",x"22",x"0A",x"26",x"22",x"65", -- 0x0980
    x"14",x"85",x"14",x"A5",x"22",x"65",x"15",x"85", -- 0x0988
    x"15",x"06",x"14",x"26",x"15",x"A5",x"14",x"65", -- 0x0990
    x"07",x"85",x"14",x"90",x"02",x"E6",x"15",x"20", -- 0x0998
    x"73",x"00",x"4C",x"71",x"C9",x"20",x"8B",x"D0", -- 0x09A0
    x"85",x"49",x"84",x"4A",x"A9",x"B2",x"20",x"FF", -- 0x09A8
    x"CE",x"A5",x"0E",x"48",x"A5",x"0D",x"48",x"20", -- 0x09B0
    x"9E",x"CD",x"68",x"2A",x"20",x"90",x"CD",x"D0", -- 0x09B8
    x"18",x"68",x"10",x"12",x"20",x"1B",x"DC",x"20", -- 0x09C0
    x"BF",x"D1",x"A0",x"00",x"A5",x"64",x"91",x"49", -- 0x09C8
    x"C8",x"A5",x"65",x"91",x"49",x"60",x"4C",x"D0", -- 0x09D0
    x"DB",x"68",x"A4",x"4A",x"C0",x"DF",x"D0",x"4C", -- 0x09D8
    x"20",x"A6",x"D6",x"C9",x"06",x"D0",x"3D",x"A0", -- 0x09E0
    x"00",x"84",x"61",x"84",x"66",x"84",x"71",x"20", -- 0x09E8
    x"1D",x"CA",x"20",x"E2",x"DA",x"E6",x"71",x"A4", -- 0x09F0
    x"71",x"20",x"1D",x"CA",x"20",x"0C",x"DC",x"AA", -- 0x09F8
    x"F0",x"05",x"E8",x"8A",x"20",x"ED",x"DA",x"A4", -- 0x0A00
    x"71",x"C8",x"C0",x"06",x"D0",x"DF",x"20",x"E2", -- 0x0A08
    x"DA",x"20",x"9B",x"DC",x"A6",x"64",x"A4",x"63", -- 0x0A10
    x"A5",x"65",x"4C",x"DB",x"FF",x"B1",x"22",x"20", -- 0x0A18
    x"80",x"00",x"90",x"03",x"4C",x"48",x"D2",x"E9", -- 0x0A20
    x"2F",x"4C",x"7E",x"DD",x"A0",x"02",x"B1",x"64", -- 0x0A28
    x"C5",x"34",x"90",x"17",x"D0",x"07",x"88",x"B1", -- 0x0A30
    x"64",x"C5",x"33",x"90",x"0E",x"A4",x"65",x"C4", -- 0x0A38
    x"2E",x"90",x"08",x"D0",x"0D",x"A5",x"64",x"C5", -- 0x0A40
    x"2D",x"B0",x"07",x"A5",x"64",x"A4",x"65",x"4C", -- 0x0A48
    x"68",x"CA",x"A0",x"00",x"B1",x"64",x"20",x"75", -- 0x0A50
    x"D4",x"A5",x"50",x"A4",x"51",x"85",x"6F",x"84", -- 0x0A58
    x"70",x"20",x"7A",x"D6",x"A9",x"61",x"A0",x"00", -- 0x0A60
    x"85",x"50",x"84",x"51",x"20",x"DB",x"D6",x"A0", -- 0x0A68
    x"00",x"B1",x"50",x"91",x"49",x"C8",x"B1",x"50", -- 0x0A70
    x"91",x"49",x"C8",x"B1",x"50",x"91",x"49",x"60", -- 0x0A78
    x"20",x"86",x"CA",x"4C",x"B5",x"CB",x"20",x"9E", -- 0x0A80
    x"D7",x"F0",x"05",x"A9",x"2C",x"20",x"FF",x"CE", -- 0x0A88
    x"08",x"86",x"13",x"20",x"15",x"E1",x"28",x"4C", -- 0x0A90
    x"A0",x"CA",x"20",x"21",x"CB",x"20",x"79",x"00", -- 0x0A98
    x"F0",x"35",x"F0",x"43",x"C9",x"A3",x"F0",x"50", -- 0x0AA0
    x"C9",x"A6",x"18",x"F0",x"4B",x"C9",x"2C",x"F0", -- 0x0AA8
    x"37",x"C9",x"3B",x"F0",x"5E",x"20",x"9E",x"CD", -- 0x0AB0
    x"24",x"0D",x"30",x"DE",x"20",x"DD",x"DD",x"20", -- 0x0AB8
    x"87",x"D4",x"20",x"21",x"CB",x"20",x"3B",x"CB", -- 0x0AC0
    x"D0",x"D3",x"A9",x"00",x"9D",x"00",x"02",x"A2", -- 0x0AC8
    x"FF",x"A0",x"01",x"A5",x"13",x"D0",x"10",x"A9", -- 0x0AD0
    x"0D",x"20",x"47",x"CB",x"24",x"13",x"10",x"05", -- 0x0AD8
    x"A9",x"0A",x"20",x"47",x"CB",x"49",x"FF",x"60", -- 0x0AE0
    x"38",x"20",x"F0",x"FF",x"98",x"38",x"E9",x"0B", -- 0x0AE8
    x"B0",x"FC",x"49",x"FF",x"69",x"01",x"D0",x"16", -- 0x0AF0
    x"08",x"38",x"20",x"F0",x"FF",x"84",x"09",x"20", -- 0x0AF8
    x"9B",x"D7",x"C9",x"29",x"D0",x"59",x"28",x"90", -- 0x0B00
    x"06",x"8A",x"E5",x"09",x"90",x"05",x"AA",x"E8", -- 0x0B08
    x"CA",x"D0",x"06",x"20",x"73",x"00",x"4C",x"A2", -- 0x0B10
    x"CA",x"20",x"3B",x"CB",x"D0",x"F2",x"20",x"87", -- 0x0B18
    x"D4",x"20",x"A6",x"D6",x"AA",x"A0",x"00",x"E8", -- 0x0B20
    x"CA",x"F0",x"BC",x"B1",x"22",x"20",x"47",x"CB", -- 0x0B28
    x"C8",x"C9",x"0D",x"D0",x"F3",x"20",x"E5",x"CA", -- 0x0B30
    x"4C",x"28",x"CB",x"A5",x"13",x"F0",x"03",x"A9", -- 0x0B38
    x"20",x"2C",x"A9",x"1D",x"2C",x"A9",x"3F",x"20", -- 0x0B40
    x"09",x"E1",x"29",x"FF",x"60",x"A5",x"11",x"F0", -- 0x0B48
    x"11",x"30",x"04",x"A0",x"FF",x"D0",x"04",x"A5", -- 0x0B50
    x"3F",x"A4",x"40",x"85",x"39",x"84",x"3A",x"4C", -- 0x0B58
    x"08",x"CF",x"A5",x"13",x"F0",x"05",x"A2",x"18", -- 0x0B60
    x"4C",x"37",x"C4",x"A9",x"0C",x"A0",x"CD",x"20", -- 0x0B68
    x"1E",x"CB",x"A5",x"3D",x"A4",x"3E",x"85",x"7A", -- 0x0B70
    x"84",x"7B",x"60",x"20",x"A6",x"D3",x"C9",x"23", -- 0x0B78
    x"D0",x"10",x"20",x"73",x"00",x"20",x"9E",x"D7", -- 0x0B80
    x"A9",x"2C",x"20",x"FF",x"CE",x"86",x"13",x"20", -- 0x0B88
    x"1B",x"E1",x"A2",x"01",x"A0",x"02",x"A9",x"00", -- 0x0B90
    x"8D",x"01",x"02",x"A9",x"40",x"20",x"0F",x"CC", -- 0x0B98
    x"A6",x"13",x"D0",x"13",x"60",x"20",x"9E",x"D7", -- 0x0BA0
    x"A9",x"2C",x"20",x"FF",x"CE",x"86",x"13",x"20", -- 0x0BA8
    x"1B",x"E1",x"20",x"CE",x"CB",x"A5",x"13",x"20", -- 0x0BB0
    x"CC",x"FF",x"A2",x"00",x"86",x"13",x"60",x"C9", -- 0x0BB8
    x"22",x"D0",x"0B",x"20",x"BD",x"CE",x"A9",x"3B", -- 0x0BC0
    x"20",x"FF",x"CE",x"20",x"21",x"CB",x"20",x"A6", -- 0x0BC8
    x"D3",x"A9",x"2C",x"8D",x"FF",x"01",x"20",x"F9", -- 0x0BD0
    x"CB",x"A5",x"13",x"F0",x"0D",x"20",x"B7",x"FF", -- 0x0BD8
    x"29",x"02",x"F0",x"06",x"20",x"B5",x"CB",x"4C", -- 0x0BE0
    x"F8",x"C8",x"AD",x"00",x"02",x"D0",x"1E",x"A5", -- 0x0BE8
    x"13",x"D0",x"E3",x"20",x"06",x"C9",x"4C",x"FB", -- 0x0BF0
    x"C8",x"A5",x"13",x"D0",x"06",x"20",x"45",x"CB", -- 0x0BF8
    x"20",x"3B",x"CB",x"4C",x"60",x"C5",x"A6",x"41", -- 0x0C00
    x"A4",x"42",x"A9",x"98",x"2C",x"A9",x"00",x"85", -- 0x0C08
    x"11",x"86",x"43",x"84",x"44",x"20",x"8B",x"D0", -- 0x0C10
    x"85",x"49",x"84",x"4A",x"A5",x"7A",x"A4",x"7B", -- 0x0C18
    x"85",x"4B",x"84",x"4C",x"A6",x"43",x"A4",x"44", -- 0x0C20
    x"86",x"7A",x"84",x"7B",x"20",x"79",x"00",x"D0", -- 0x0C28
    x"20",x"24",x"11",x"50",x"0C",x"20",x"21",x"E1", -- 0x0C30
    x"8D",x"00",x"02",x"A2",x"FF",x"A0",x"01",x"D0", -- 0x0C38
    x"0C",x"30",x"75",x"A5",x"13",x"D0",x"03",x"20", -- 0x0C40
    x"45",x"CB",x"20",x"F9",x"CB",x"86",x"7A",x"84", -- 0x0C48
    x"7B",x"20",x"73",x"00",x"24",x"0D",x"10",x"31", -- 0x0C50
    x"24",x"11",x"50",x"09",x"E8",x"86",x"7A",x"A9", -- 0x0C58
    x"00",x"85",x"07",x"F0",x"0C",x"85",x"07",x"C9", -- 0x0C60
    x"22",x"F0",x"07",x"A9",x"3A",x"85",x"07",x"A9", -- 0x0C68
    x"2C",x"18",x"85",x"08",x"A5",x"7A",x"A4",x"7B", -- 0x0C70
    x"69",x"00",x"90",x"01",x"C8",x"20",x"8D",x"D4", -- 0x0C78
    x"20",x"E2",x"D7",x"20",x"DA",x"C9",x"4C",x"91", -- 0x0C80
    x"CC",x"20",x"F3",x"DC",x"A5",x"0E",x"20",x"C2", -- 0x0C88
    x"C9",x"20",x"79",x"00",x"F0",x"07",x"C9",x"2C", -- 0x0C90
    x"F0",x"03",x"4C",x"4D",x"CB",x"A5",x"7A",x"A4", -- 0x0C98
    x"7B",x"85",x"43",x"84",x"44",x"A5",x"4B",x"A4", -- 0x0CA0
    x"4C",x"85",x"7A",x"84",x"7B",x"20",x"79",x"00", -- 0x0CA8
    x"F0",x"2D",x"20",x"FD",x"CE",x"4C",x"15",x"CC", -- 0x0CB0
    x"20",x"06",x"C9",x"C8",x"AA",x"D0",x"12",x"A2", -- 0x0CB8
    x"0D",x"C8",x"B1",x"7A",x"F0",x"6C",x"C8",x"B1", -- 0x0CC0
    x"7A",x"85",x"3F",x"C8",x"B1",x"7A",x"C8",x"85", -- 0x0CC8
    x"40",x"20",x"FB",x"C8",x"20",x"79",x"00",x"AA", -- 0x0CD0
    x"E0",x"83",x"D0",x"DC",x"4C",x"51",x"CC",x"A5", -- 0x0CD8
    x"43",x"A4",x"44",x"A6",x"11",x"10",x"03",x"4C", -- 0x0CE0
    x"27",x"C8",x"A0",x"00",x"B1",x"43",x"F0",x"0B", -- 0x0CE8
    x"A5",x"13",x"D0",x"07",x"A9",x"FC",x"A0",x"CC", -- 0x0CF0
    x"4C",x"1E",x"CB",x"60",x"3F",x"45",x"58",x"54", -- 0x0CF8
    x"52",x"41",x"20",x"49",x"47",x"4E",x"4F",x"52", -- 0x0D00
    x"45",x"44",x"0D",x"00",x"3F",x"52",x"45",x"44", -- 0x0D08
    x"4F",x"20",x"46",x"52",x"4F",x"4D",x"20",x"53", -- 0x0D10
    x"54",x"41",x"52",x"54",x"0D",x"00",x"D0",x"04", -- 0x0D18
    x"A0",x"00",x"F0",x"03",x"20",x"8B",x"D0",x"85", -- 0x0D20
    x"49",x"84",x"4A",x"20",x"8A",x"C3",x"F0",x"05", -- 0x0D28
    x"A2",x"0A",x"4C",x"37",x"C4",x"9A",x"8A",x"18", -- 0x0D30
    x"69",x"04",x"48",x"69",x"06",x"85",x"24",x"68", -- 0x0D38
    x"A0",x"01",x"20",x"A2",x"DB",x"BA",x"BD",x"09", -- 0x0D40
    x"01",x"85",x"66",x"A5",x"49",x"A4",x"4A",x"20", -- 0x0D48
    x"67",x"D8",x"20",x"D0",x"DB",x"A0",x"01",x"20", -- 0x0D50
    x"5D",x"DC",x"BA",x"38",x"FD",x"09",x"01",x"F0", -- 0x0D58
    x"17",x"BD",x"0F",x"01",x"85",x"39",x"BD",x"10", -- 0x0D60
    x"01",x"85",x"3A",x"BD",x"12",x"01",x"85",x"7A", -- 0x0D68
    x"BD",x"11",x"01",x"85",x"7B",x"4C",x"AE",x"C7", -- 0x0D70
    x"8A",x"69",x"11",x"AA",x"9A",x"20",x"79",x"00", -- 0x0D78
    x"C9",x"2C",x"D0",x"F1",x"20",x"73",x"00",x"20", -- 0x0D80
    x"24",x"CD",x"20",x"9E",x"CD",x"18",x"24",x"38", -- 0x0D88
    x"24",x"0D",x"30",x"03",x"B0",x"03",x"60",x"B0", -- 0x0D90
    x"FD",x"A2",x"16",x"4C",x"37",x"C4",x"A6",x"7A", -- 0x0D98
    x"D0",x"02",x"C6",x"7B",x"C6",x"7A",x"A2",x"00", -- 0x0DA0
    x"24",x"48",x"8A",x"48",x"A9",x"01",x"20",x"FB", -- 0x0DA8
    x"C3",x"20",x"83",x"CE",x"A9",x"00",x"85",x"4D", -- 0x0DB0
    x"20",x"79",x"00",x"38",x"E9",x"B1",x"90",x"17", -- 0x0DB8
    x"C9",x"03",x"B0",x"13",x"C9",x"01",x"2A",x"49", -- 0x0DC0
    x"01",x"45",x"4D",x"C5",x"4D",x"90",x"61",x"85", -- 0x0DC8
    x"4D",x"20",x"73",x"00",x"4C",x"BB",x"CD",x"A6", -- 0x0DD0
    x"4D",x"D0",x"2C",x"B0",x"7B",x"69",x"07",x"90", -- 0x0DD8
    x"77",x"65",x"0D",x"D0",x"03",x"4C",x"3D",x"D6", -- 0x0DE0
    x"69",x"FF",x"85",x"22",x"0A",x"65",x"22",x"A8", -- 0x0DE8
    x"68",x"D9",x"80",x"C0",x"B0",x"67",x"20",x"8D", -- 0x0DF0
    x"CD",x"48",x"20",x"20",x"CE",x"68",x"A4",x"4B", -- 0x0DF8
    x"10",x"17",x"AA",x"F0",x"56",x"D0",x"5F",x"46", -- 0x0E00
    x"0D",x"8A",x"2A",x"A6",x"7A",x"D0",x"02",x"C6", -- 0x0E08
    x"7B",x"C6",x"7A",x"A0",x"1B",x"85",x"4D",x"D0", -- 0x0E10
    x"D7",x"D9",x"80",x"C0",x"B0",x"48",x"90",x"D9", -- 0x0E18
    x"B9",x"82",x"C0",x"48",x"B9",x"81",x"C0",x"48", -- 0x0E20
    x"20",x"33",x"CE",x"A5",x"4D",x"4C",x"A9",x"CD", -- 0x0E28
    x"4C",x"08",x"CF",x"A5",x"66",x"BE",x"80",x"C0", -- 0x0E30
    x"A8",x"68",x"85",x"22",x"E6",x"22",x"68",x"85", -- 0x0E38
    x"23",x"98",x"48",x"20",x"1B",x"DC",x"A5",x"65", -- 0x0E40
    x"48",x"A5",x"64",x"48",x"A5",x"63",x"48",x"A5", -- 0x0E48
    x"62",x"48",x"A5",x"61",x"48",x"6C",x"22",x"00", -- 0x0E50
    x"A0",x"FF",x"68",x"F0",x"23",x"C9",x"64",x"F0", -- 0x0E58
    x"03",x"20",x"8D",x"CD",x"84",x"4B",x"68",x"4A", -- 0x0E60
    x"85",x"12",x"68",x"85",x"69",x"68",x"85",x"6A", -- 0x0E68
    x"68",x"85",x"6B",x"68",x"85",x"6C",x"68",x"85", -- 0x0E70
    x"6D",x"68",x"85",x"6E",x"45",x"66",x"85",x"6F", -- 0x0E78
    x"A5",x"61",x"60",x"6C",x"0A",x"03",x"A9",x"00", -- 0x0E80
    x"85",x"0D",x"20",x"73",x"00",x"B0",x"03",x"4C", -- 0x0E88
    x"F3",x"DC",x"20",x"13",x"D1",x"90",x"03",x"4C", -- 0x0E90
    x"28",x"CF",x"C9",x"FF",x"D0",x"0F",x"A9",x"A8", -- 0x0E98
    x"A0",x"CE",x"20",x"A2",x"DB",x"4C",x"73",x"00", -- 0x0EA0
    x"82",x"49",x"0F",x"DA",x"A1",x"C9",x"2E",x"F0", -- 0x0EA8
    x"DE",x"C9",x"AB",x"F0",x"58",x"C9",x"AA",x"F0", -- 0x0EB0
    x"D1",x"C9",x"22",x"D0",x"0F",x"A5",x"7A",x"A4", -- 0x0EB8
    x"7B",x"69",x"00",x"90",x"01",x"C8",x"20",x"87", -- 0x0EC0
    x"D4",x"4C",x"E2",x"D7",x"C9",x"A8",x"D0",x"13", -- 0x0EC8
    x"A0",x"18",x"D0",x"3B",x"20",x"BF",x"D1",x"A5", -- 0x0ED0
    x"65",x"49",x"FF",x"A8",x"A5",x"64",x"49",x"FF", -- 0x0ED8
    x"4C",x"91",x"D3",x"C9",x"A5",x"D0",x"03",x"4C", -- 0x0EE0
    x"F4",x"D3",x"C9",x"B4",x"90",x"03",x"4C",x"A7", -- 0x0EE8
    x"CF",x"20",x"FA",x"CE",x"20",x"9E",x"CD",x"A9", -- 0x0EF0
    x"29",x"2C",x"A9",x"28",x"2C",x"A9",x"2C",x"A0", -- 0x0EF8
    x"00",x"D1",x"7A",x"D0",x"03",x"4C",x"73",x"00", -- 0x0F00
    x"A2",x"0B",x"4C",x"37",x"C4",x"A0",x"15",x"68", -- 0x0F08
    x"68",x"4C",x"FA",x"CD",x"38",x"A5",x"64",x"E9", -- 0x0F10
    x"00",x"A5",x"65",x"E9",x"C0",x"90",x"08",x"A9", -- 0x0F18
    x"87",x"E5",x"64",x"A9",x"E3",x"E5",x"65",x"60", -- 0x0F20
    x"20",x"8B",x"D0",x"85",x"64",x"84",x"65",x"A6", -- 0x0F28
    x"45",x"A4",x"46",x"A5",x"0D",x"F0",x"26",x"A9", -- 0x0F30
    x"00",x"85",x"70",x"20",x"14",x"CF",x"90",x"1C", -- 0x0F38
    x"E0",x"54",x"D0",x"18",x"C0",x"C9",x"D0",x"14", -- 0x0F40
    x"20",x"84",x"CF",x"84",x"5E",x"88",x"84",x"71", -- 0x0F48
    x"A0",x"06",x"84",x"5D",x"A0",x"24",x"20",x"68", -- 0x0F50
    x"DE",x"4C",x"6F",x"D4",x"60",x"24",x"0E",x"10", -- 0x0F58
    x"0D",x"A0",x"00",x"B1",x"64",x"AA",x"C8",x"B1", -- 0x0F60
    x"64",x"A8",x"8A",x"4C",x"91",x"D3",x"20",x"14", -- 0x0F68
    x"CF",x"90",x"2D",x"E0",x"54",x"D0",x"1B",x"C0", -- 0x0F70
    x"49",x"D0",x"25",x"20",x"84",x"CF",x"98",x"A2", -- 0x0F78
    x"A0",x"4C",x"4F",x"DC",x"20",x"DE",x"FF",x"86", -- 0x0F80
    x"64",x"84",x"63",x"85",x"65",x"A0",x"00",x"84", -- 0x0F88
    x"62",x"60",x"E0",x"53",x"D0",x"0A",x"C0",x"54", -- 0x0F90
    x"D0",x"06",x"20",x"B7",x"FF",x"4C",x"3C",x"DC", -- 0x0F98
    x"A5",x"64",x"A4",x"65",x"4C",x"A2",x"DB",x"0A", -- 0x0FA0
    x"48",x"AA",x"20",x"73",x"00",x"E0",x"8F",x"90", -- 0x0FA8
    x"20",x"20",x"FA",x"CE",x"20",x"9E",x"CD",x"20", -- 0x0FB0
    x"FD",x"CE",x"20",x"8F",x"CD",x"68",x"AA",x"A5", -- 0x0FB8
    x"65",x"48",x"A5",x"64",x"48",x"8A",x"48",x"20", -- 0x0FC0
    x"9E",x"D7",x"68",x"A8",x"8A",x"48",x"4C",x"D6", -- 0x0FC8
    x"CF",x"20",x"F1",x"CE",x"68",x"A8",x"B9",x"EA", -- 0x0FD0
    x"BF",x"85",x"55",x"B9",x"EB",x"BF",x"85",x"56", -- 0x0FD8
    x"20",x"54",x"00",x"4C",x"8D",x"CD",x"A0",x"FF", -- 0x0FE0
    x"2C",x"A0",x"00",x"84",x"0B",x"20",x"BF",x"D1", -- 0x0FE8
    x"A5",x"64",x"45",x"0B",x"85",x"07",x"A5",x"65", -- 0x0FF0
    x"45",x"0B",x"85",x"08",x"20",x"FC",x"DB",x"20", -- 0x0FF8
    x"BF",x"D1",x"A5",x"65",x"45",x"0B",x"25",x"08", -- 0x1000
    x"45",x"0B",x"A8",x"A5",x"64",x"45",x"0B",x"25", -- 0x1008
    x"07",x"45",x"0B",x"4C",x"91",x"D3",x"20",x"90", -- 0x1010
    x"CD",x"B0",x"13",x"A5",x"6E",x"09",x"7F",x"25", -- 0x1018
    x"6A",x"85",x"6A",x"A9",x"69",x"A0",x"00",x"20", -- 0x1020
    x"5B",x"DC",x"AA",x"4C",x"61",x"D0",x"A9",x"00", -- 0x1028
    x"85",x"0D",x"C6",x"4D",x"20",x"A6",x"D6",x"85", -- 0x1030
    x"61",x"86",x"62",x"84",x"63",x"A5",x"6C",x"A4", -- 0x1038
    x"6D",x"20",x"AA",x"D6",x"86",x"6C",x"84",x"6D", -- 0x1040
    x"AA",x"38",x"E5",x"61",x"F0",x"08",x"A9",x"01", -- 0x1048
    x"90",x"04",x"A6",x"61",x"A9",x"FF",x"85",x"66", -- 0x1050
    x"A0",x"FF",x"E8",x"C8",x"CA",x"D0",x"07",x"A6", -- 0x1058
    x"66",x"30",x"0F",x"18",x"90",x"0C",x"B1",x"6C", -- 0x1060
    x"D1",x"62",x"F0",x"EF",x"A2",x"FF",x"B0",x"02", -- 0x1068
    x"A2",x"01",x"E8",x"8A",x"2A",x"25",x"12",x"F0", -- 0x1070
    x"02",x"A9",x"FF",x"4C",x"3C",x"DC",x"20",x"FD", -- 0x1078
    x"CE",x"AA",x"20",x"90",x"D0",x"20",x"79",x"00", -- 0x1080
    x"D0",x"F4",x"60",x"A2",x"00",x"20",x"79",x"00", -- 0x1088
    x"86",x"0C",x"85",x"45",x"20",x"79",x"00",x"20", -- 0x1090
    x"13",x"D1",x"B0",x"03",x"4C",x"08",x"CF",x"A2", -- 0x1098
    x"00",x"86",x"0D",x"86",x"0E",x"20",x"73",x"00", -- 0x10A0
    x"90",x"05",x"20",x"13",x"D1",x"90",x"0B",x"AA", -- 0x10A8
    x"20",x"73",x"00",x"90",x"FB",x"20",x"13",x"D1", -- 0x10B0
    x"B0",x"F6",x"C9",x"24",x"D0",x"06",x"A9",x"FF", -- 0x10B8
    x"85",x"0D",x"D0",x"10",x"C9",x"25",x"D0",x"13", -- 0x10C0
    x"A5",x"10",x"D0",x"D0",x"A9",x"80",x"85",x"0E", -- 0x10C8
    x"05",x"45",x"85",x"45",x"8A",x"09",x"80",x"AA", -- 0x10D0
    x"20",x"73",x"00",x"86",x"46",x"38",x"05",x"10", -- 0x10D8
    x"E9",x"28",x"D0",x"03",x"4C",x"D1",x"D1",x"A0", -- 0x10E0
    x"00",x"84",x"10",x"A5",x"2D",x"A6",x"2E",x"86", -- 0x10E8
    x"60",x"85",x"5F",x"E4",x"30",x"D0",x"04",x"C5", -- 0x10F0
    x"2F",x"F0",x"22",x"A5",x"45",x"D1",x"5F",x"D0", -- 0x10F8
    x"08",x"A5",x"46",x"C8",x"D1",x"5F",x"F0",x"7D", -- 0x1100
    x"88",x"18",x"A5",x"5F",x"69",x"07",x"90",x"E1", -- 0x1108
    x"E8",x"D0",x"DC",x"C9",x"41",x"90",x"05",x"E9", -- 0x1110
    x"5B",x"38",x"E9",x"A5",x"60",x"68",x"48",x"C9", -- 0x1118
    x"2A",x"D0",x"05",x"A9",x"13",x"A0",x"DF",x"60", -- 0x1120
    x"A5",x"45",x"A4",x"46",x"C9",x"54",x"D0",x"0B", -- 0x1128
    x"C0",x"C9",x"F0",x"EF",x"C0",x"49",x"D0",x"03", -- 0x1130
    x"4C",x"08",x"CF",x"C9",x"53",x"D0",x"04",x"C0", -- 0x1138
    x"54",x"F0",x"F5",x"A5",x"2F",x"A4",x"30",x"85", -- 0x1140
    x"5F",x"84",x"60",x"A5",x"31",x"A4",x"32",x"85", -- 0x1148
    x"5A",x"84",x"5B",x"18",x"69",x"07",x"90",x"01", -- 0x1150
    x"C8",x"85",x"58",x"84",x"59",x"20",x"B8",x"C3", -- 0x1158
    x"A5",x"58",x"A4",x"59",x"C8",x"85",x"2F",x"84", -- 0x1160
    x"30",x"A0",x"00",x"A5",x"45",x"91",x"5F",x"C8", -- 0x1168
    x"A5",x"46",x"91",x"5F",x"A9",x"00",x"C8",x"91", -- 0x1170
    x"5F",x"C8",x"91",x"5F",x"C8",x"91",x"5F",x"C8", -- 0x1178
    x"91",x"5F",x"C8",x"91",x"5F",x"A5",x"5F",x"18", -- 0x1180
    x"69",x"02",x"A4",x"60",x"90",x"01",x"C8",x"85", -- 0x1188
    x"47",x"84",x"48",x"60",x"A5",x"0B",x"0A",x"69", -- 0x1190
    x"05",x"65",x"5F",x"A4",x"60",x"90",x"01",x"C8", -- 0x1198
    x"85",x"58",x"84",x"59",x"60",x"90",x"80",x"00", -- 0x11A0
    x"00",x"00",x"20",x"BF",x"D1",x"A5",x"64",x"A4", -- 0x11A8
    x"65",x"60",x"20",x"73",x"00",x"20",x"9E",x"CD", -- 0x11B0
    x"20",x"8D",x"CD",x"A5",x"66",x"30",x"0D",x"A5", -- 0x11B8
    x"61",x"C9",x"90",x"90",x"09",x"A9",x"A5",x"A0", -- 0x11C0
    x"D1",x"20",x"5B",x"DC",x"D0",x"7A",x"4C",x"9B", -- 0x11C8
    x"DC",x"A5",x"0C",x"05",x"0E",x"48",x"A5",x"0D", -- 0x11D0
    x"48",x"A0",x"00",x"98",x"48",x"A5",x"46",x"48", -- 0x11D8
    x"A5",x"45",x"48",x"20",x"B2",x"D1",x"68",x"85", -- 0x11E0
    x"45",x"68",x"85",x"46",x"68",x"A8",x"BA",x"BD", -- 0x11E8
    x"02",x"01",x"48",x"BD",x"01",x"01",x"48",x"A5", -- 0x11F0
    x"64",x"9D",x"02",x"01",x"A5",x"65",x"9D",x"01", -- 0x11F8
    x"01",x"C8",x"20",x"79",x"00",x"C9",x"2C",x"F0", -- 0x1200
    x"D2",x"84",x"0B",x"20",x"F7",x"CE",x"68",x"85", -- 0x1208
    x"0D",x"68",x"85",x"0E",x"29",x"7F",x"85",x"0C", -- 0x1210
    x"A6",x"2F",x"A5",x"30",x"86",x"5F",x"85",x"60", -- 0x1218
    x"C5",x"32",x"D0",x"04",x"E4",x"31",x"F0",x"39", -- 0x1220
    x"A0",x"00",x"B1",x"5F",x"C8",x"C5",x"45",x"D0", -- 0x1228
    x"06",x"A5",x"46",x"D1",x"5F",x"F0",x"16",x"C8", -- 0x1230
    x"B1",x"5F",x"18",x"65",x"5F",x"AA",x"C8",x"B1", -- 0x1238
    x"5F",x"65",x"60",x"90",x"D7",x"A2",x"12",x"2C", -- 0x1240
    x"A2",x"0E",x"4C",x"37",x"C4",x"A2",x"13",x"A5", -- 0x1248
    x"0C",x"D0",x"F7",x"20",x"94",x"D1",x"A5",x"0B", -- 0x1250
    x"A0",x"04",x"D1",x"5F",x"D0",x"E7",x"4C",x"EA", -- 0x1258
    x"D2",x"20",x"94",x"D1",x"20",x"08",x"C4",x"A0", -- 0x1260
    x"00",x"84",x"72",x"A2",x"05",x"A5",x"45",x"91", -- 0x1268
    x"5F",x"10",x"01",x"CA",x"C8",x"A5",x"46",x"91", -- 0x1270
    x"5F",x"10",x"02",x"CA",x"CA",x"86",x"71",x"A5", -- 0x1278
    x"0B",x"C8",x"C8",x"C8",x"91",x"5F",x"A2",x"0B", -- 0x1280
    x"A9",x"00",x"24",x"0C",x"50",x"08",x"68",x"18", -- 0x1288
    x"69",x"01",x"AA",x"68",x"69",x"00",x"C8",x"91", -- 0x1290
    x"5F",x"C8",x"8A",x"91",x"5F",x"20",x"4C",x"D3", -- 0x1298
    x"86",x"71",x"85",x"72",x"A4",x"22",x"C6",x"0B", -- 0x12A0
    x"D0",x"DC",x"65",x"59",x"B0",x"5D",x"85",x"59", -- 0x12A8
    x"A8",x"8A",x"65",x"58",x"90",x"03",x"C8",x"F0", -- 0x12B0
    x"52",x"20",x"08",x"C4",x"85",x"31",x"84",x"32", -- 0x12B8
    x"A9",x"00",x"E6",x"72",x"A4",x"71",x"F0",x"05", -- 0x12C0
    x"88",x"91",x"58",x"D0",x"FB",x"C6",x"59",x"C6", -- 0x12C8
    x"72",x"D0",x"F5",x"E6",x"59",x"38",x"A5",x"31", -- 0x12D0
    x"E5",x"5F",x"A0",x"02",x"91",x"5F",x"A5",x"32", -- 0x12D8
    x"C8",x"E5",x"60",x"91",x"5F",x"A5",x"0C",x"D0", -- 0x12E0
    x"62",x"C8",x"B1",x"5F",x"85",x"0B",x"A9",x"00", -- 0x12E8
    x"85",x"71",x"85",x"72",x"C8",x"68",x"AA",x"85", -- 0x12F0
    x"64",x"68",x"85",x"65",x"D1",x"5F",x"90",x"0E", -- 0x12F8
    x"D0",x"06",x"C8",x"8A",x"D1",x"5F",x"90",x"07", -- 0x1300
    x"4C",x"45",x"D2",x"4C",x"35",x"C4",x"C8",x"A5", -- 0x1308
    x"72",x"05",x"71",x"18",x"F0",x"0A",x"20",x"4C", -- 0x1310
    x"D3",x"8A",x"65",x"64",x"AA",x"98",x"A4",x"22", -- 0x1318
    x"65",x"65",x"86",x"71",x"C6",x"0B",x"D0",x"CA", -- 0x1320
    x"85",x"72",x"A2",x"05",x"A5",x"45",x"10",x"01", -- 0x1328
    x"CA",x"A5",x"46",x"10",x"02",x"CA",x"CA",x"86", -- 0x1330
    x"28",x"A9",x"00",x"20",x"55",x"D3",x"8A",x"65", -- 0x1338
    x"58",x"85",x"47",x"98",x"65",x"59",x"85",x"48", -- 0x1340
    x"A8",x"A5",x"47",x"60",x"84",x"22",x"B1",x"5F", -- 0x1348
    x"85",x"28",x"88",x"B1",x"5F",x"85",x"29",x"A9", -- 0x1350
    x"10",x"85",x"5D",x"A2",x"00",x"A0",x"00",x"8A", -- 0x1358
    x"0A",x"AA",x"98",x"2A",x"A8",x"B0",x"A4",x"06", -- 0x1360
    x"71",x"26",x"72",x"90",x"0B",x"18",x"8A",x"65", -- 0x1368
    x"28",x"AA",x"98",x"65",x"29",x"A8",x"B0",x"93", -- 0x1370
    x"C6",x"5D",x"D0",x"E3",x"60",x"A5",x"0D",x"F0", -- 0x1378
    x"03",x"20",x"A6",x"D6",x"20",x"26",x"D5",x"38", -- 0x1380
    x"A5",x"33",x"E5",x"31",x"A8",x"A5",x"34",x"E5", -- 0x1388
    x"32",x"A2",x"00",x"86",x"0D",x"85",x"62",x"84", -- 0x1390
    x"63",x"A2",x"90",x"4C",x"44",x"DC",x"38",x"20", -- 0x1398
    x"F0",x"FF",x"A9",x"00",x"F0",x"EB",x"A6",x"3A", -- 0x13A0
    x"E8",x"D0",x"A0",x"A2",x"15",x"2C",x"A2",x"1B", -- 0x13A8
    x"4C",x"37",x"C4",x"20",x"E1",x"D3",x"20",x"A6", -- 0x13B0
    x"D3",x"20",x"FA",x"CE",x"A9",x"80",x"85",x"10", -- 0x13B8
    x"20",x"8B",x"D0",x"20",x"8D",x"CD",x"20",x"F7", -- 0x13C0
    x"CE",x"A9",x"B2",x"20",x"FF",x"CE",x"48",x"A5", -- 0x13C8
    x"48",x"48",x"A5",x"47",x"48",x"A5",x"7B",x"48", -- 0x13D0
    x"A5",x"7A",x"48",x"20",x"F8",x"C8",x"4C",x"4F", -- 0x13D8
    x"D4",x"A9",x"A5",x"20",x"FF",x"CE",x"09",x"80", -- 0x13E0
    x"85",x"10",x"20",x"92",x"D0",x"85",x"4E",x"84", -- 0x13E8
    x"4F",x"4C",x"8D",x"CD",x"20",x"E1",x"D3",x"A5", -- 0x13F0
    x"4F",x"48",x"A5",x"4E",x"48",x"20",x"F1",x"CE", -- 0x13F8
    x"20",x"8D",x"CD",x"68",x"85",x"4E",x"68",x"85", -- 0x1400
    x"4F",x"A0",x"02",x"B1",x"4E",x"85",x"47",x"AA", -- 0x1408
    x"C8",x"B1",x"4E",x"F0",x"99",x"85",x"48",x"C8", -- 0x1410
    x"B1",x"47",x"48",x"88",x"10",x"FA",x"A4",x"48", -- 0x1418
    x"20",x"D4",x"DB",x"A5",x"7B",x"48",x"A5",x"7A", -- 0x1420
    x"48",x"B1",x"4E",x"85",x"7A",x"C8",x"B1",x"4E", -- 0x1428
    x"85",x"7B",x"A5",x"48",x"48",x"A5",x"47",x"48", -- 0x1430
    x"20",x"8A",x"CD",x"68",x"85",x"4E",x"68",x"85", -- 0x1438
    x"4F",x"20",x"79",x"00",x"F0",x"03",x"4C",x"08", -- 0x1440
    x"CF",x"68",x"85",x"7A",x"68",x"85",x"7B",x"A0", -- 0x1448
    x"00",x"68",x"91",x"4E",x"68",x"C8",x"91",x"4E", -- 0x1450
    x"68",x"C8",x"91",x"4E",x"68",x"C8",x"91",x"4E", -- 0x1458
    x"68",x"C8",x"91",x"4E",x"60",x"20",x"8D",x"CD", -- 0x1460
    x"A0",x"00",x"20",x"DF",x"DD",x"68",x"68",x"A9", -- 0x1468
    x"FF",x"A0",x"00",x"F0",x"12",x"A6",x"64",x"A4", -- 0x1470
    x"65",x"86",x"50",x"84",x"51",x"20",x"F4",x"D4", -- 0x1478
    x"86",x"62",x"84",x"63",x"85",x"61",x"60",x"A2", -- 0x1480
    x"22",x"86",x"07",x"86",x"08",x"85",x"6F",x"84", -- 0x1488
    x"70",x"85",x"62",x"84",x"63",x"A0",x"FF",x"C8", -- 0x1490
    x"B1",x"6F",x"F0",x"0C",x"C5",x"07",x"F0",x"04", -- 0x1498
    x"C5",x"08",x"D0",x"F3",x"C9",x"22",x"F0",x"01", -- 0x14A0
    x"18",x"84",x"61",x"98",x"65",x"6F",x"85",x"71", -- 0x14A8
    x"A6",x"70",x"90",x"01",x"E8",x"86",x"72",x"A5", -- 0x14B0
    x"70",x"F0",x"04",x"C9",x"02",x"D0",x"0B",x"98", -- 0x14B8
    x"20",x"75",x"D4",x"A6",x"6F",x"A4",x"70",x"20", -- 0x14C0
    x"88",x"D6",x"A6",x"16",x"E0",x"22",x"D0",x"05", -- 0x14C8
    x"A2",x"19",x"4C",x"37",x"C4",x"A5",x"61",x"95", -- 0x14D0
    x"00",x"A5",x"62",x"95",x"01",x"A5",x"63",x"95", -- 0x14D8
    x"02",x"A0",x"00",x"86",x"64",x"84",x"65",x"84", -- 0x14E0
    x"70",x"88",x"84",x"0D",x"86",x"17",x"E8",x"E8", -- 0x14E8
    x"E8",x"86",x"16",x"60",x"46",x"0F",x"48",x"49", -- 0x14F0
    x"FF",x"38",x"65",x"33",x"A4",x"34",x"B0",x"01", -- 0x14F8
    x"88",x"C4",x"32",x"90",x"11",x"D0",x"04",x"C5", -- 0x1500
    x"31",x"90",x"0B",x"85",x"33",x"84",x"34",x"85", -- 0x1508
    x"35",x"84",x"36",x"AA",x"68",x"60",x"A2",x"10", -- 0x1510
    x"A5",x"0F",x"30",x"B6",x"20",x"26",x"D5",x"A9", -- 0x1518
    x"80",x"85",x"0F",x"68",x"D0",x"D0",x"A6",x"37", -- 0x1520
    x"A5",x"38",x"86",x"33",x"85",x"34",x"A0",x"00", -- 0x1528
    x"84",x"4F",x"84",x"4E",x"A5",x"31",x"A6",x"32", -- 0x1530
    x"85",x"5F",x"86",x"60",x"A9",x"19",x"A2",x"00", -- 0x1538
    x"85",x"22",x"86",x"23",x"C5",x"16",x"F0",x"05", -- 0x1540
    x"20",x"C7",x"D5",x"F0",x"F7",x"A9",x"07",x"85", -- 0x1548
    x"53",x"A5",x"2D",x"A6",x"2E",x"85",x"22",x"86", -- 0x1550
    x"23",x"E4",x"30",x"D0",x"04",x"C5",x"2F",x"F0", -- 0x1558
    x"05",x"20",x"BD",x"D5",x"F0",x"F3",x"85",x"58", -- 0x1560
    x"86",x"59",x"A9",x"03",x"85",x"53",x"A5",x"58", -- 0x1568
    x"A6",x"59",x"E4",x"32",x"D0",x"07",x"C5",x"31", -- 0x1570
    x"D0",x"03",x"4C",x"06",x"D6",x"85",x"22",x"86", -- 0x1578
    x"23",x"A0",x"00",x"B1",x"22",x"AA",x"C8",x"B1", -- 0x1580
    x"22",x"08",x"C8",x"B1",x"22",x"65",x"58",x"85", -- 0x1588
    x"58",x"C8",x"B1",x"22",x"65",x"59",x"85",x"59", -- 0x1590
    x"28",x"10",x"D3",x"8A",x"30",x"D0",x"C8",x"B1", -- 0x1598
    x"22",x"A0",x"00",x"0A",x"69",x"05",x"65",x"22", -- 0x15A0
    x"85",x"22",x"90",x"02",x"E6",x"23",x"A6",x"23", -- 0x15A8
    x"E4",x"59",x"D0",x"04",x"C5",x"58",x"F0",x"BA", -- 0x15B0
    x"20",x"C7",x"D5",x"F0",x"F3",x"B1",x"22",x"30", -- 0x15B8
    x"35",x"C8",x"B1",x"22",x"10",x"30",x"C8",x"B1", -- 0x15C0
    x"22",x"F0",x"2B",x"C8",x"B1",x"22",x"AA",x"C8", -- 0x15C8
    x"B1",x"22",x"C5",x"34",x"90",x"06",x"D0",x"1E", -- 0x15D0
    x"E4",x"33",x"B0",x"1A",x"C5",x"60",x"90",x"16", -- 0x15D8
    x"D0",x"04",x"E4",x"5F",x"90",x"10",x"86",x"5F", -- 0x15E0
    x"85",x"60",x"A5",x"22",x"A6",x"23",x"85",x"4E", -- 0x15E8
    x"86",x"4F",x"A5",x"53",x"85",x"55",x"A5",x"53", -- 0x15F0
    x"18",x"65",x"22",x"85",x"22",x"90",x"02",x"E6", -- 0x15F8
    x"23",x"A6",x"23",x"A0",x"00",x"60",x"A5",x"4F", -- 0x1600
    x"05",x"4E",x"F0",x"F5",x"A5",x"55",x"29",x"04", -- 0x1608
    x"4A",x"A8",x"85",x"55",x"B1",x"4E",x"65",x"5F", -- 0x1610
    x"85",x"5A",x"A5",x"60",x"69",x"00",x"85",x"5B", -- 0x1618
    x"A5",x"33",x"A6",x"34",x"85",x"58",x"86",x"59", -- 0x1620
    x"20",x"BF",x"C3",x"A4",x"55",x"C8",x"A5",x"58", -- 0x1628
    x"91",x"4E",x"AA",x"E6",x"59",x"A5",x"59",x"C8", -- 0x1630
    x"91",x"4E",x"4C",x"2A",x"D5",x"A5",x"65",x"48", -- 0x1638
    x"A5",x"64",x"48",x"20",x"83",x"CE",x"20",x"8F", -- 0x1640
    x"CD",x"68",x"85",x"6F",x"68",x"85",x"70",x"A0", -- 0x1648
    x"00",x"B1",x"6F",x"18",x"71",x"64",x"90",x"05", -- 0x1650
    x"A2",x"17",x"4C",x"37",x"C4",x"20",x"75",x"D4", -- 0x1658
    x"20",x"7A",x"D6",x"A5",x"50",x"A4",x"51",x"20", -- 0x1660
    x"AA",x"D6",x"20",x"8C",x"D6",x"A5",x"6F",x"A4", -- 0x1668
    x"70",x"20",x"AA",x"D6",x"20",x"CA",x"D4",x"4C", -- 0x1670
    x"B8",x"CD",x"A0",x"00",x"B1",x"6F",x"48",x"C8", -- 0x1678
    x"B1",x"6F",x"AA",x"C8",x"B1",x"6F",x"A8",x"68", -- 0x1680
    x"86",x"22",x"84",x"23",x"A8",x"F0",x"0A",x"48", -- 0x1688
    x"88",x"B1",x"22",x"91",x"35",x"98",x"D0",x"F8", -- 0x1690
    x"68",x"18",x"65",x"35",x"85",x"35",x"90",x"02", -- 0x1698
    x"E6",x"36",x"60",x"20",x"8F",x"CD",x"A5",x"64", -- 0x16A0
    x"A4",x"65",x"85",x"22",x"84",x"23",x"20",x"DB", -- 0x16A8
    x"D6",x"08",x"A0",x"00",x"B1",x"22",x"48",x"C8", -- 0x16B0
    x"B1",x"22",x"AA",x"C8",x"B1",x"22",x"A8",x"68", -- 0x16B8
    x"28",x"D0",x"13",x"C4",x"34",x"D0",x"0F",x"E4", -- 0x16C0
    x"33",x"D0",x"0B",x"48",x"18",x"65",x"33",x"85", -- 0x16C8
    x"33",x"90",x"02",x"E6",x"34",x"68",x"86",x"22", -- 0x16D0
    x"84",x"23",x"60",x"C4",x"18",x"D0",x"0C",x"C5", -- 0x16D8
    x"17",x"D0",x"08",x"85",x"16",x"E9",x"03",x"85", -- 0x16E0
    x"17",x"A0",x"00",x"60",x"20",x"A1",x"D7",x"8A", -- 0x16E8
    x"48",x"A9",x"01",x"20",x"7D",x"D4",x"68",x"A0", -- 0x16F0
    x"00",x"91",x"62",x"68",x"68",x"4C",x"CA",x"D4", -- 0x16F8
    x"20",x"61",x"D7",x"D1",x"50",x"98",x"90",x"04", -- 0x1700
    x"B1",x"50",x"AA",x"98",x"48",x"8A",x"48",x"20", -- 0x1708
    x"7D",x"D4",x"A5",x"50",x"A4",x"51",x"20",x"AA", -- 0x1710
    x"D6",x"68",x"A8",x"68",x"18",x"65",x"22",x"85", -- 0x1718
    x"22",x"90",x"02",x"E6",x"23",x"98",x"20",x"8C", -- 0x1720
    x"D6",x"4C",x"CA",x"D4",x"20",x"61",x"D7",x"18", -- 0x1728
    x"F1",x"50",x"49",x"FF",x"4C",x"06",x"D7",x"A9", -- 0x1730
    x"FF",x"85",x"65",x"20",x"79",x"00",x"C9",x"29", -- 0x1738
    x"F0",x"06",x"20",x"FD",x"CE",x"20",x"9E",x"D7", -- 0x1740
    x"20",x"61",x"D7",x"F0",x"4B",x"CA",x"8A",x"48", -- 0x1748
    x"18",x"A2",x"00",x"F1",x"50",x"B0",x"B6",x"49", -- 0x1750
    x"FF",x"C5",x"65",x"90",x"B1",x"A5",x"65",x"B0", -- 0x1758
    x"AD",x"20",x"F7",x"CE",x"68",x"A8",x"68",x"85", -- 0x1760
    x"55",x"68",x"68",x"68",x"AA",x"68",x"85",x"50", -- 0x1768
    x"68",x"85",x"51",x"A5",x"55",x"48",x"98",x"48", -- 0x1770
    x"A0",x"00",x"8A",x"60",x"20",x"82",x"D7",x"4C", -- 0x1778
    x"A2",x"D3",x"20",x"A3",x"D6",x"A2",x"00",x"86", -- 0x1780
    x"0D",x"A8",x"60",x"20",x"82",x"D7",x"F0",x"08", -- 0x1788
    x"A0",x"00",x"B1",x"22",x"A8",x"4C",x"A2",x"D3", -- 0x1790
    x"4C",x"48",x"D2",x"20",x"73",x"00",x"20",x"8A", -- 0x1798
    x"CD",x"20",x"B8",x"D1",x"A6",x"64",x"D0",x"F0", -- 0x17A0
    x"A6",x"65",x"4C",x"79",x"00",x"20",x"82",x"D7", -- 0x17A8
    x"D0",x"03",x"4C",x"F7",x"D8",x"A6",x"7A",x"A4", -- 0x17B0
    x"7B",x"86",x"71",x"84",x"72",x"A6",x"22",x"86", -- 0x17B8
    x"7A",x"18",x"65",x"22",x"85",x"24",x"A6",x"23", -- 0x17C0
    x"86",x"7B",x"90",x"01",x"E8",x"86",x"25",x"A0", -- 0x17C8
    x"00",x"B1",x"24",x"48",x"98",x"91",x"24",x"20", -- 0x17D0
    x"79",x"00",x"20",x"F3",x"DC",x"68",x"A0",x"00", -- 0x17D8
    x"91",x"24",x"A6",x"71",x"A4",x"72",x"86",x"7A", -- 0x17E0
    x"84",x"7B",x"60",x"20",x"8A",x"CD",x"20",x"F7", -- 0x17E8
    x"D7",x"20",x"FD",x"CE",x"4C",x"9E",x"D7",x"A5", -- 0x17F0
    x"66",x"30",x"9D",x"A5",x"61",x"C9",x"91",x"B0", -- 0x17F8
    x"97",x"20",x"9B",x"DC",x"A5",x"64",x"A4",x"65", -- 0x1800
    x"84",x"14",x"85",x"15",x"60",x"A5",x"15",x"48", -- 0x1808
    x"A5",x"14",x"48",x"20",x"F7",x"D7",x"A0",x"00", -- 0x1810
    x"B1",x"14",x"A8",x"68",x"85",x"14",x"68",x"85", -- 0x1818
    x"15",x"4C",x"A2",x"D3",x"20",x"EB",x"D7",x"8A", -- 0x1820
    x"A0",x"00",x"91",x"14",x"60",x"20",x"EB",x"D7", -- 0x1828
    x"86",x"49",x"A2",x"00",x"20",x"79",x"00",x"F0", -- 0x1830
    x"03",x"20",x"F1",x"D7",x"86",x"4A",x"A0",x"00", -- 0x1838
    x"B1",x"14",x"45",x"4A",x"25",x"49",x"F0",x"F8", -- 0x1840
    x"60",x"A9",x"11",x"A0",x"DF",x"4C",x"67",x"D8", -- 0x1848
    x"20",x"8C",x"DA",x"A5",x"66",x"49",x"FF",x"85", -- 0x1850
    x"66",x"45",x"6E",x"85",x"6F",x"A5",x"61",x"4C", -- 0x1858
    x"6A",x"D8",x"20",x"99",x"D9",x"90",x"3C",x"20", -- 0x1860
    x"8C",x"DA",x"D0",x"03",x"4C",x"FC",x"DB",x"A6", -- 0x1868
    x"70",x"86",x"56",x"A2",x"69",x"A5",x"69",x"A8", -- 0x1870
    x"F0",x"CE",x"38",x"E5",x"61",x"F0",x"24",x"90", -- 0x1878
    x"12",x"84",x"61",x"A4",x"6E",x"84",x"66",x"49", -- 0x1880
    x"FF",x"69",x"00",x"A0",x"00",x"84",x"56",x"A2", -- 0x1888
    x"61",x"D0",x"04",x"A0",x"00",x"84",x"70",x"C9", -- 0x1890
    x"F9",x"30",x"C7",x"A8",x"A5",x"70",x"56",x"01", -- 0x1898
    x"20",x"B0",x"D9",x"24",x"6F",x"10",x"57",x"A0", -- 0x18A0
    x"61",x"E0",x"69",x"F0",x"02",x"A0",x"69",x"38", -- 0x18A8
    x"49",x"FF",x"65",x"56",x"85",x"70",x"B9",x"04", -- 0x18B0
    x"00",x"F5",x"04",x"85",x"65",x"B9",x"03",x"00", -- 0x18B8
    x"F5",x"03",x"85",x"64",x"B9",x"02",x"00",x"F5", -- 0x18C0
    x"02",x"85",x"63",x"B9",x"01",x"00",x"F5",x"01", -- 0x18C8
    x"85",x"62",x"B0",x"03",x"20",x"47",x"D9",x"A0", -- 0x18D0
    x"00",x"98",x"18",x"A6",x"62",x"D0",x"4A",x"A6", -- 0x18D8
    x"63",x"86",x"62",x"A6",x"64",x"86",x"63",x"A6", -- 0x18E0
    x"65",x"86",x"64",x"A6",x"70",x"86",x"65",x"84", -- 0x18E8
    x"70",x"69",x"08",x"C9",x"20",x"D0",x"E4",x"A9", -- 0x18F0
    x"00",x"85",x"61",x"85",x"66",x"60",x"65",x"56", -- 0x18F8
    x"85",x"70",x"A5",x"65",x"65",x"6D",x"85",x"65", -- 0x1900
    x"A5",x"64",x"65",x"6C",x"85",x"64",x"A5",x"63", -- 0x1908
    x"65",x"6B",x"85",x"63",x"A5",x"62",x"65",x"6A", -- 0x1910
    x"85",x"62",x"4C",x"36",x"D9",x"69",x"01",x"06", -- 0x1918
    x"70",x"26",x"65",x"26",x"64",x"26",x"63",x"26", -- 0x1920
    x"62",x"10",x"F2",x"38",x"E5",x"61",x"B0",x"C7", -- 0x1928
    x"49",x"FF",x"69",x"01",x"85",x"61",x"90",x"0E", -- 0x1930
    x"E6",x"61",x"F0",x"42",x"66",x"62",x"66",x"63", -- 0x1938
    x"66",x"64",x"66",x"65",x"66",x"70",x"60",x"A5", -- 0x1940
    x"66",x"49",x"FF",x"85",x"66",x"A5",x"62",x"49", -- 0x1948
    x"FF",x"85",x"62",x"A5",x"63",x"49",x"FF",x"85", -- 0x1950
    x"63",x"A5",x"64",x"49",x"FF",x"85",x"64",x"A5", -- 0x1958
    x"65",x"49",x"FF",x"85",x"65",x"A5",x"70",x"49", -- 0x1960
    x"FF",x"85",x"70",x"E6",x"70",x"D0",x"0E",x"E6", -- 0x1968
    x"65",x"D0",x"0A",x"E6",x"64",x"D0",x"06",x"E6", -- 0x1970
    x"63",x"D0",x"02",x"E6",x"62",x"60",x"A2",x"0F", -- 0x1978
    x"4C",x"37",x"C4",x"A2",x"25",x"B4",x"04",x"84", -- 0x1980
    x"70",x"B4",x"03",x"94",x"04",x"B4",x"02",x"94", -- 0x1988
    x"03",x"B4",x"01",x"94",x"02",x"A4",x"68",x"94", -- 0x1990
    x"01",x"69",x"08",x"30",x"E8",x"F0",x"E6",x"E9", -- 0x1998
    x"08",x"A8",x"A5",x"70",x"B0",x"14",x"16",x"01", -- 0x19A0
    x"90",x"02",x"F6",x"01",x"76",x"01",x"76",x"01", -- 0x19A8
    x"76",x"02",x"76",x"03",x"76",x"04",x"6A",x"C8", -- 0x19B0
    x"D0",x"EC",x"18",x"60",x"81",x"00",x"00",x"00", -- 0x19B8
    x"00",x"03",x"7F",x"5E",x"56",x"CB",x"79",x"80", -- 0x19C0
    x"13",x"9B",x"0B",x"64",x"80",x"76",x"38",x"93", -- 0x19C8
    x"16",x"82",x"38",x"AA",x"3B",x"20",x"80",x"35", -- 0x19D0
    x"04",x"F3",x"34",x"81",x"35",x"04",x"F3",x"34", -- 0x19D8
    x"80",x"80",x"00",x"00",x"00",x"80",x"31",x"72", -- 0x19E0
    x"17",x"F8",x"20",x"2B",x"DC",x"F0",x"02",x"10", -- 0x19E8
    x"03",x"4C",x"48",x"D2",x"A5",x"61",x"E9",x"7F", -- 0x19F0
    x"48",x"A9",x"80",x"85",x"61",x"A9",x"D6",x"A0", -- 0x19F8
    x"D9",x"20",x"67",x"D8",x"A9",x"DB",x"A0",x"D9", -- 0x1A00
    x"20",x"0F",x"DB",x"A9",x"BC",x"A0",x"D9",x"20", -- 0x1A08
    x"50",x"D8",x"A9",x"C1",x"A0",x"D9",x"20",x"40", -- 0x1A10
    x"E0",x"A9",x"E0",x"A0",x"D9",x"20",x"67",x"D8", -- 0x1A18
    x"68",x"20",x"7E",x"DD",x"A9",x"E5",x"A0",x"D9", -- 0x1A20
    x"20",x"8C",x"DA",x"D0",x"03",x"4C",x"8B",x"DA", -- 0x1A28
    x"20",x"B7",x"DA",x"A9",x"00",x"85",x"26",x"85", -- 0x1A30
    x"27",x"85",x"28",x"85",x"29",x"A5",x"70",x"20", -- 0x1A38
    x"59",x"DA",x"A5",x"65",x"20",x"59",x"DA",x"A5", -- 0x1A40
    x"64",x"20",x"59",x"DA",x"A5",x"63",x"20",x"59", -- 0x1A48
    x"DA",x"A5",x"62",x"20",x"5E",x"DA",x"4C",x"8F", -- 0x1A50
    x"DB",x"D0",x"03",x"4C",x"83",x"D9",x"4A",x"09", -- 0x1A58
    x"80",x"A8",x"90",x"19",x"18",x"A5",x"29",x"65", -- 0x1A60
    x"6D",x"85",x"29",x"A5",x"28",x"65",x"6C",x"85", -- 0x1A68
    x"28",x"A5",x"27",x"65",x"6B",x"85",x"27",x"A5", -- 0x1A70
    x"26",x"65",x"6A",x"85",x"26",x"66",x"26",x"66", -- 0x1A78
    x"27",x"66",x"28",x"66",x"29",x"66",x"70",x"98", -- 0x1A80
    x"4A",x"D0",x"D6",x"60",x"85",x"22",x"84",x"23", -- 0x1A88
    x"A0",x"04",x"B1",x"22",x"85",x"6D",x"88",x"B1", -- 0x1A90
    x"22",x"85",x"6C",x"88",x"B1",x"22",x"85",x"6B", -- 0x1A98
    x"88",x"B1",x"22",x"85",x"6E",x"45",x"66",x"85", -- 0x1AA0
    x"6F",x"A5",x"6E",x"09",x"80",x"85",x"6A",x"88", -- 0x1AA8
    x"B1",x"22",x"85",x"69",x"A5",x"61",x"60",x"A5", -- 0x1AB0
    x"69",x"F0",x"1F",x"18",x"65",x"61",x"90",x"04", -- 0x1AB8
    x"30",x"1D",x"18",x"2C",x"10",x"14",x"69",x"80", -- 0x1AC0
    x"85",x"61",x"D0",x"03",x"4C",x"FB",x"D8",x"A5", -- 0x1AC8
    x"6F",x"85",x"66",x"60",x"A5",x"66",x"49",x"FF", -- 0x1AD0
    x"30",x"05",x"68",x"68",x"4C",x"F7",x"D8",x"4C", -- 0x1AD8
    x"7E",x"D9",x"20",x"0C",x"DC",x"AA",x"F0",x"10", -- 0x1AE0
    x"18",x"69",x"02",x"B0",x"F2",x"A2",x"00",x"86", -- 0x1AE8
    x"6F",x"20",x"77",x"D8",x"E6",x"61",x"F0",x"E7", -- 0x1AF0
    x"60",x"84",x"20",x"00",x"00",x"00",x"20",x"0C", -- 0x1AF8
    x"DC",x"A9",x"F9",x"A0",x"DA",x"A2",x"00",x"86", -- 0x1B00
    x"6F",x"20",x"A2",x"DB",x"4C",x"12",x"DB",x"20", -- 0x1B08
    x"8C",x"DA",x"F0",x"76",x"20",x"1B",x"DC",x"A9", -- 0x1B10
    x"00",x"38",x"E5",x"61",x"85",x"61",x"20",x"B7", -- 0x1B18
    x"DA",x"E6",x"61",x"F0",x"BA",x"A2",x"FC",x"A9", -- 0x1B20
    x"01",x"A4",x"6A",x"C4",x"62",x"D0",x"10",x"A4", -- 0x1B28
    x"6B",x"C4",x"63",x"D0",x"0A",x"A4",x"6C",x"C4", -- 0x1B30
    x"64",x"D0",x"04",x"A4",x"6D",x"C4",x"65",x"08", -- 0x1B38
    x"2A",x"90",x"09",x"E8",x"95",x"29",x"F0",x"32", -- 0x1B40
    x"10",x"34",x"A9",x"01",x"28",x"B0",x"0E",x"06", -- 0x1B48
    x"6D",x"26",x"6C",x"26",x"6B",x"26",x"6A",x"B0", -- 0x1B50
    x"E6",x"30",x"CE",x"10",x"E2",x"A8",x"A5",x"6D", -- 0x1B58
    x"E5",x"65",x"85",x"6D",x"A5",x"6C",x"E5",x"64", -- 0x1B60
    x"85",x"6C",x"A5",x"6B",x"E5",x"63",x"85",x"6B", -- 0x1B68
    x"A5",x"6A",x"E5",x"62",x"85",x"6A",x"98",x"4C", -- 0x1B70
    x"4F",x"DB",x"A9",x"40",x"D0",x"CE",x"0A",x"0A", -- 0x1B78
    x"0A",x"0A",x"0A",x"0A",x"85",x"70",x"28",x"4C", -- 0x1B80
    x"8F",x"DB",x"A2",x"14",x"4C",x"37",x"C4",x"A5", -- 0x1B88
    x"26",x"85",x"62",x"A5",x"27",x"85",x"63",x"A5", -- 0x1B90
    x"28",x"85",x"64",x"A5",x"29",x"85",x"65",x"4C", -- 0x1B98
    x"D7",x"D8",x"85",x"22",x"84",x"23",x"A0",x"04", -- 0x1BA0
    x"B1",x"22",x"85",x"65",x"88",x"B1",x"22",x"85", -- 0x1BA8
    x"64",x"88",x"B1",x"22",x"85",x"63",x"88",x"B1", -- 0x1BB0
    x"22",x"85",x"66",x"09",x"80",x"85",x"62",x"88", -- 0x1BB8
    x"B1",x"22",x"85",x"61",x"84",x"70",x"60",x"A2", -- 0x1BC0
    x"5C",x"2C",x"A2",x"57",x"A0",x"00",x"F0",x"04", -- 0x1BC8
    x"A6",x"49",x"A4",x"4A",x"20",x"1B",x"DC",x"86", -- 0x1BD0
    x"22",x"84",x"23",x"A0",x"04",x"A5",x"65",x"91", -- 0x1BD8
    x"22",x"88",x"A5",x"64",x"91",x"22",x"88",x"A5", -- 0x1BE0
    x"63",x"91",x"22",x"88",x"A5",x"66",x"09",x"7F", -- 0x1BE8
    x"25",x"62",x"91",x"22",x"88",x"A5",x"61",x"91", -- 0x1BF0
    x"22",x"84",x"70",x"60",x"A5",x"6E",x"85",x"66", -- 0x1BF8
    x"A2",x"05",x"B5",x"68",x"95",x"60",x"CA",x"D0", -- 0x1C00
    x"F9",x"86",x"70",x"60",x"20",x"1B",x"DC",x"A2", -- 0x1C08
    x"06",x"B5",x"60",x"95",x"68",x"CA",x"D0",x"F9", -- 0x1C10
    x"86",x"70",x"60",x"A5",x"61",x"F0",x"FB",x"06", -- 0x1C18
    x"70",x"90",x"F7",x"20",x"6F",x"D9",x"D0",x"F2", -- 0x1C20
    x"4C",x"38",x"D9",x"A5",x"61",x"F0",x"09",x"A5", -- 0x1C28
    x"66",x"2A",x"A9",x"FF",x"B0",x"02",x"A9",x"01", -- 0x1C30
    x"60",x"20",x"2B",x"DC",x"85",x"62",x"A9",x"00", -- 0x1C38
    x"85",x"63",x"A2",x"88",x"A5",x"62",x"49",x"FF", -- 0x1C40
    x"2A",x"A9",x"00",x"85",x"65",x"85",x"64",x"86", -- 0x1C48
    x"61",x"85",x"70",x"85",x"66",x"4C",x"D2",x"D8", -- 0x1C50
    x"46",x"66",x"60",x"85",x"24",x"84",x"25",x"A0", -- 0x1C58
    x"00",x"B1",x"24",x"C8",x"AA",x"F0",x"C4",x"B1", -- 0x1C60
    x"24",x"45",x"66",x"30",x"C2",x"E4",x"61",x"D0", -- 0x1C68
    x"21",x"B1",x"24",x"09",x"80",x"C5",x"62",x"D0", -- 0x1C70
    x"19",x"C8",x"B1",x"24",x"C5",x"63",x"D0",x"12", -- 0x1C78
    x"C8",x"B1",x"24",x"C5",x"64",x"D0",x"0B",x"C8", -- 0x1C80
    x"A9",x"7F",x"C5",x"70",x"B1",x"24",x"E5",x"65", -- 0x1C88
    x"F0",x"28",x"A5",x"66",x"90",x"02",x"49",x"FF", -- 0x1C90
    x"4C",x"31",x"DC",x"A5",x"61",x"F0",x"4A",x"38", -- 0x1C98
    x"E9",x"A0",x"24",x"66",x"10",x"09",x"AA",x"A9", -- 0x1CA0
    x"FF",x"85",x"68",x"20",x"4D",x"D9",x"8A",x"A2", -- 0x1CA8
    x"61",x"C9",x"F9",x"10",x"06",x"20",x"99",x"D9", -- 0x1CB0
    x"84",x"68",x"60",x"A8",x"A5",x"66",x"29",x"80", -- 0x1CB8
    x"46",x"62",x"05",x"62",x"85",x"62",x"20",x"B0", -- 0x1CC0
    x"D9",x"84",x"68",x"60",x"A5",x"61",x"C9",x"A0", -- 0x1CC8
    x"B0",x"20",x"20",x"9B",x"DC",x"84",x"70",x"A5", -- 0x1CD0
    x"66",x"84",x"66",x"49",x"80",x"2A",x"A9",x"A0", -- 0x1CD8
    x"85",x"61",x"A5",x"65",x"85",x"07",x"4C",x"D2", -- 0x1CE0
    x"D8",x"85",x"62",x"85",x"63",x"85",x"64",x"85", -- 0x1CE8
    x"65",x"A8",x"60",x"A0",x"00",x"A2",x"0A",x"94", -- 0x1CF0
    x"5D",x"CA",x"10",x"FB",x"90",x"0F",x"C9",x"2D", -- 0x1CF8
    x"D0",x"04",x"86",x"67",x"F0",x"04",x"C9",x"2B", -- 0x1D00
    x"D0",x"05",x"20",x"73",x"00",x"90",x"5B",x"C9", -- 0x1D08
    x"2E",x"F0",x"2E",x"C9",x"45",x"D0",x"30",x"20", -- 0x1D10
    x"73",x"00",x"90",x"17",x"C9",x"AB",x"F0",x"0E", -- 0x1D18
    x"C9",x"2D",x"F0",x"0A",x"C9",x"AA",x"F0",x"08", -- 0x1D20
    x"C9",x"2B",x"F0",x"04",x"D0",x"07",x"66",x"60", -- 0x1D28
    x"20",x"73",x"00",x"90",x"5C",x"24",x"60",x"10", -- 0x1D30
    x"0E",x"A9",x"00",x"38",x"E5",x"5E",x"4C",x"49", -- 0x1D38
    x"DD",x"66",x"5F",x"24",x"5F",x"50",x"C3",x"A5", -- 0x1D40
    x"5E",x"38",x"E5",x"5D",x"85",x"5E",x"F0",x"12", -- 0x1D48
    x"10",x"09",x"20",x"FE",x"DA",x"E6",x"5E",x"D0", -- 0x1D50
    x"F9",x"F0",x"07",x"20",x"E2",x"DA",x"C6",x"5E", -- 0x1D58
    x"D0",x"F9",x"A5",x"67",x"30",x"01",x"60",x"4C", -- 0x1D60
    x"B4",x"DF",x"48",x"24",x"5F",x"10",x"02",x"E6", -- 0x1D68
    x"5D",x"20",x"E2",x"DA",x"68",x"38",x"E9",x"30", -- 0x1D70
    x"20",x"7E",x"DD",x"4C",x"0A",x"DD",x"48",x"20", -- 0x1D78
    x"0C",x"DC",x"68",x"20",x"3C",x"DC",x"A5",x"6E", -- 0x1D80
    x"45",x"66",x"85",x"6F",x"A6",x"61",x"4C",x"6A", -- 0x1D88
    x"D8",x"A5",x"5E",x"C9",x"0A",x"90",x"09",x"A9", -- 0x1D90
    x"64",x"24",x"60",x"30",x"11",x"4C",x"7E",x"D9", -- 0x1D98
    x"0A",x"0A",x"18",x"65",x"5E",x"0A",x"18",x"A0", -- 0x1DA0
    x"00",x"71",x"7A",x"38",x"E9",x"30",x"85",x"5E", -- 0x1DA8
    x"4C",x"30",x"DD",x"9B",x"3E",x"BC",x"1F",x"FD", -- 0x1DB0
    x"9E",x"6E",x"6B",x"27",x"FD",x"9E",x"6E",x"6B", -- 0x1DB8
    x"28",x"00",x"A9",x"71",x"A0",x"C3",x"20",x"DA", -- 0x1DC0
    x"DD",x"A5",x"3A",x"A6",x"39",x"85",x"62",x"86", -- 0x1DC8
    x"63",x"A2",x"90",x"38",x"20",x"49",x"DC",x"20", -- 0x1DD0
    x"DF",x"DD",x"4C",x"1E",x"CB",x"A0",x"01",x"A9", -- 0x1DD8
    x"20",x"24",x"66",x"10",x"02",x"A9",x"2D",x"99", -- 0x1DE0
    x"FF",x"00",x"85",x"66",x"84",x"71",x"C8",x"A9", -- 0x1DE8
    x"30",x"A6",x"61",x"D0",x"03",x"4C",x"04",x"DF", -- 0x1DF0
    x"A9",x"00",x"E0",x"80",x"F0",x"02",x"B0",x"09", -- 0x1DF8
    x"A9",x"BD",x"A0",x"DD",x"20",x"28",x"DA",x"A9", -- 0x1E00
    x"F7",x"85",x"5D",x"A9",x"B8",x"A0",x"DD",x"20", -- 0x1E08
    x"5B",x"DC",x"F0",x"1E",x"10",x"12",x"A9",x"B3", -- 0x1E10
    x"A0",x"DD",x"20",x"5B",x"DC",x"F0",x"02",x"10", -- 0x1E18
    x"0E",x"20",x"E2",x"DA",x"C6",x"5D",x"D0",x"EE", -- 0x1E20
    x"20",x"FE",x"DA",x"E6",x"5D",x"D0",x"DC",x"20", -- 0x1E28
    x"49",x"D8",x"20",x"9B",x"DC",x"A2",x"01",x"A5", -- 0x1E30
    x"5D",x"18",x"69",x"0A",x"30",x"09",x"C9",x"0B", -- 0x1E38
    x"B0",x"06",x"69",x"FF",x"AA",x"A9",x"02",x"38", -- 0x1E40
    x"E9",x"02",x"85",x"5E",x"86",x"5D",x"8A",x"F0", -- 0x1E48
    x"02",x"10",x"13",x"A4",x"71",x"A9",x"2E",x"C8", -- 0x1E50
    x"99",x"FF",x"00",x"8A",x"F0",x"06",x"A9",x"30", -- 0x1E58
    x"C8",x"99",x"FF",x"00",x"84",x"71",x"A0",x"00", -- 0x1E60
    x"A2",x"80",x"A5",x"65",x"18",x"79",x"19",x"DF", -- 0x1E68
    x"85",x"65",x"A5",x"64",x"79",x"18",x"DF",x"85", -- 0x1E70
    x"64",x"A5",x"63",x"79",x"17",x"DF",x"85",x"63", -- 0x1E78
    x"A5",x"62",x"79",x"16",x"DF",x"85",x"62",x"E8", -- 0x1E80
    x"B0",x"04",x"10",x"DE",x"30",x"02",x"30",x"DA", -- 0x1E88
    x"8A",x"90",x"04",x"49",x"FF",x"69",x"0A",x"69", -- 0x1E90
    x"2F",x"C8",x"C8",x"C8",x"C8",x"84",x"47",x"A4", -- 0x1E98
    x"71",x"C8",x"AA",x"29",x"7F",x"99",x"FF",x"00", -- 0x1EA0
    x"C6",x"5D",x"D0",x"06",x"A9",x"2E",x"C8",x"99", -- 0x1EA8
    x"FF",x"00",x"84",x"71",x"A4",x"47",x"8A",x"49", -- 0x1EB0
    x"FF",x"29",x"80",x"AA",x"C0",x"24",x"F0",x"04", -- 0x1EB8
    x"C0",x"3C",x"D0",x"A6",x"A4",x"71",x"B9",x"FF", -- 0x1EC0
    x"00",x"88",x"C9",x"30",x"F0",x"F8",x"C9",x"2E", -- 0x1EC8
    x"F0",x"01",x"C8",x"A9",x"2B",x"A6",x"5E",x"F0", -- 0x1ED0
    x"2E",x"10",x"08",x"A9",x"00",x"38",x"E5",x"5E", -- 0x1ED8
    x"AA",x"A9",x"2D",x"99",x"01",x"01",x"A9",x"45", -- 0x1EE0
    x"99",x"00",x"01",x"8A",x"A2",x"2F",x"38",x"E8", -- 0x1EE8
    x"E9",x"0A",x"B0",x"FB",x"69",x"3A",x"99",x"03", -- 0x1EF0
    x"01",x"8A",x"99",x"02",x"01",x"A9",x"00",x"99", -- 0x1EF8
    x"04",x"01",x"F0",x"08",x"99",x"FF",x"00",x"A9", -- 0x1F00
    x"00",x"99",x"00",x"01",x"A9",x"00",x"A0",x"01", -- 0x1F08
    x"60",x"80",x"00",x"00",x"00",x"00",x"FA",x"0A", -- 0x1F10
    x"1F",x"00",x"00",x"98",x"96",x"80",x"FF",x"F0", -- 0x1F18
    x"BD",x"C0",x"00",x"01",x"86",x"A0",x"FF",x"FF", -- 0x1F20
    x"D8",x"F0",x"00",x"00",x"03",x"E8",x"FF",x"FF", -- 0x1F28
    x"FF",x"9C",x"00",x"00",x"00",x"0A",x"FF",x"FF", -- 0x1F30
    x"FF",x"FF",x"FF",x"DF",x"0A",x"80",x"00",x"03", -- 0x1F38
    x"4B",x"C0",x"FF",x"FF",x"73",x"60",x"00",x"00", -- 0x1F40
    x"0E",x"10",x"FF",x"FF",x"FD",x"A8",x"00",x"00", -- 0x1F48
    x"00",x"3C",x"BF",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x1F50
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x1F58
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x1F60
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x1F68
    x"AA",x"20",x"0C",x"DC",x"A9",x"11",x"A0",x"DF", -- 0x1F70
    x"20",x"A2",x"DB",x"F0",x"70",x"A5",x"69",x"D0", -- 0x1F78
    x"03",x"4C",x"F9",x"D8",x"A2",x"4E",x"A0",x"00", -- 0x1F80
    x"20",x"D4",x"DB",x"A5",x"6E",x"10",x"0F",x"20", -- 0x1F88
    x"CC",x"DC",x"A9",x"4E",x"A0",x"00",x"20",x"5B", -- 0x1F90
    x"DC",x"D0",x"03",x"98",x"A4",x"07",x"20",x"FE", -- 0x1F98
    x"DB",x"98",x"48",x"20",x"EA",x"D9",x"A9",x"4E", -- 0x1FA0
    x"A0",x"00",x"20",x"28",x"DA",x"20",x"ED",x"DF", -- 0x1FA8
    x"68",x"4A",x"90",x"0A",x"A5",x"61",x"F0",x"06", -- 0x1FB0
    x"A5",x"66",x"49",x"FF",x"85",x"66",x"60",x"81", -- 0x1FB8
    x"38",x"AA",x"3B",x"29",x"07",x"71",x"34",x"58", -- 0x1FC0
    x"3E",x"56",x"74",x"16",x"7E",x"B3",x"1B",x"77", -- 0x1FC8
    x"2F",x"EE",x"E3",x"85",x"7A",x"1D",x"84",x"1C", -- 0x1FD0
    x"2A",x"7C",x"63",x"59",x"58",x"0A",x"7E",x"75", -- 0x1FD8
    x"FD",x"E7",x"C6",x"80",x"31",x"72",x"18",x"10", -- 0x1FE0
    x"81",x"00",x"00",x"00",x"00",x"A9",x"BF",x"A0", -- 0x1FE8
    x"DF",x"20",x"28",x"DA",x"A5",x"70",x"69",x"50", -- 0x1FF0
    x"90",x"03",x"20",x"23",x"DC",x"85",x"56",x"20"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
