-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_PGM_45 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_PGM_45 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"3A",x"18",x"81",x"A7",x"C8",x"11",x"06",x"A8", -- 0x0000
    x"06",x"08",x"21",x"9C",x"24",x"7E",x"12",x"23", -- 0x0008
    x"13",x"7E",x"12",x"23",x"C5",x"01",x"1F",x"00", -- 0x0010
    x"EB",x"09",x"EB",x"C1",x"10",x"EF",x"AF",x"32", -- 0x0018
    x"18",x"81",x"C9",x"2A",x"00",x"80",x"01",x"32", -- 0x0020
    x"20",x"26",x"00",x"29",x"09",x"4E",x"23",x"66", -- 0x0028
    x"69",x"E9",x"48",x"20",x"E1",x"20",x"04",x"21", -- 0x0030
    x"24",x"21",x"44",x"21",x"64",x"21",x"81",x"21", -- 0x0038
    x"A1",x"21",x"C1",x"21",x"E1",x"21",x"01",x"22", -- 0x0040
    x"21",x"70",x"82",x"7E",x"23",x"46",x"23",x"4E", -- 0x0048
    x"2A",x"76",x"24",x"11",x"8C",x"24",x"DD",x"21", -- 0x0050
    x"00",x"81",x"FD",x"21",x"00",x"81",x"32",x"B1", -- 0x0058
    x"81",x"ED",x"53",x"01",x"80",x"E5",x"C5",x"D5", -- 0x0060
    x"CD",x"21",x"22",x"3A",x"5B",x"82",x"A7",x"20", -- 0x0068
    x"0B",x"79",x"2F",x"3C",x"DD",x"77",x"01",x"DD", -- 0x0070
    x"23",x"FD",x"34",x"00",x"D1",x"C1",x"E1",x"78", -- 0x0078
    x"32",x"03",x"80",x"1A",x"77",x"23",x"13",x"1A", -- 0x0080
    x"77",x"2B",x"D5",x"11",x"20",x"00",x"19",x"D1", -- 0x0088
    x"10",x"1A",x"3A",x"B1",x"81",x"5F",x"16",x"00", -- 0x0090
    x"19",x"0D",x"C2",x"B0",x"20",x"21",x"00",x"80", -- 0x0098
    x"34",x"7E",x"FE",x"0B",x"DA",x"23",x"20",x"AF", -- 0x00A0
    x"77",x"C3",x"BB",x"20",x"13",x"C3",x"83",x"20", -- 0x00A8
    x"ED",x"5B",x"01",x"80",x"3A",x"03",x"80",x"47", -- 0x00B0
    x"C3",x"65",x"20",x"C9",x"01",x"FF",x"03",x"21", -- 0x00B8
    x"00",x"A8",x"3A",x"00",x"88",x"36",x"28",x"23", -- 0x00C0
    x"0B",x"78",x"A7",x"20",x"F5",x"79",x"A7",x"20", -- 0x00C8
    x"F1",x"01",x"FF",x"EF",x"3A",x"00",x"88",x"0B", -- 0x00D0
    x"78",x"A7",x"20",x"F8",x"79",x"A7",x"20",x"F4", -- 0x00D8
    x"C9",x"CD",x"00",x"20",x"21",x"73",x"82",x"7E", -- 0x00E0
    x"23",x"46",x"23",x"4E",x"2A",x"78",x"24",x"11", -- 0x00E8
    x"AC",x"24",x"DD",x"21",x"09",x"81",x"FD",x"21", -- 0x00F0
    x"09",x"81",x"32",x"B1",x"81",x"ED",x"53",x"01", -- 0x00F8
    x"80",x"C3",x"65",x"20",x"21",x"76",x"82",x"7E", -- 0x0100
    x"23",x"46",x"23",x"4E",x"2A",x"7A",x"24",x"11", -- 0x0108
    x"C4",x"24",x"DD",x"21",x"12",x"81",x"FD",x"21", -- 0x0110
    x"12",x"81",x"32",x"B1",x"81",x"ED",x"53",x"01", -- 0x0118
    x"80",x"C3",x"65",x"20",x"21",x"79",x"82",x"7E", -- 0x0120
    x"23",x"46",x"23",x"4E",x"2A",x"7C",x"24",x"11", -- 0x0128
    x"DC",x"24",x"DD",x"21",x"1B",x"81",x"FD",x"21", -- 0x0130
    x"1B",x"81",x"32",x"B1",x"81",x"ED",x"53",x"01", -- 0x0138
    x"80",x"C3",x"65",x"20",x"21",x"7C",x"82",x"7E", -- 0x0140
    x"23",x"46",x"23",x"4E",x"2A",x"7E",x"24",x"11", -- 0x0148
    x"E8",x"24",x"DD",x"21",x"24",x"81",x"FD",x"21", -- 0x0150
    x"24",x"81",x"32",x"B1",x"81",x"ED",x"53",x"01", -- 0x0158
    x"80",x"C3",x"65",x"20",x"C3",x"9D",x"20",x"11", -- 0x0160
    x"24",x"25",x"01",x"04",x"02",x"DD",x"21",x"2D", -- 0x0168
    x"81",x"FD",x"21",x"2D",x"81",x"3E",x"80",x"32", -- 0x0170
    x"B1",x"81",x"ED",x"53",x"01",x"80",x"C3",x"65", -- 0x0178
    x"20",x"21",x"82",x"82",x"7E",x"23",x"46",x"23", -- 0x0180
    x"4E",x"2A",x"82",x"24",x"11",x"28",x"25",x"DD", -- 0x0188
    x"21",x"36",x"81",x"FD",x"21",x"36",x"81",x"32", -- 0x0190
    x"B1",x"81",x"ED",x"53",x"01",x"80",x"C3",x"65", -- 0x0198
    x"20",x"21",x"85",x"82",x"7E",x"23",x"46",x"23", -- 0x01A0
    x"4E",x"2A",x"84",x"24",x"11",x"30",x"25",x"DD", -- 0x01A8
    x"21",x"3F",x"81",x"FD",x"21",x"3F",x"81",x"32", -- 0x01B0
    x"B1",x"81",x"ED",x"53",x"01",x"80",x"C3",x"65", -- 0x01B8
    x"20",x"21",x"88",x"82",x"7E",x"23",x"46",x"23", -- 0x01C0
    x"4E",x"2A",x"86",x"24",x"11",x"34",x"25",x"DD", -- 0x01C8
    x"21",x"48",x"81",x"FD",x"21",x"48",x"81",x"32", -- 0x01D0
    x"B1",x"81",x"ED",x"53",x"01",x"80",x"C3",x"65", -- 0x01D8
    x"20",x"21",x"8B",x"82",x"7E",x"23",x"46",x"23", -- 0x01E0
    x"4E",x"2A",x"88",x"24",x"11",x"38",x"25",x"DD", -- 0x01E8
    x"21",x"51",x"81",x"FD",x"21",x"51",x"81",x"32", -- 0x01F0
    x"B1",x"81",x"ED",x"53",x"01",x"80",x"C3",x"65", -- 0x01F8
    x"20",x"21",x"8E",x"82",x"7E",x"23",x"46",x"23", -- 0x0200
    x"4E",x"2A",x"8A",x"24",x"11",x"3C",x"25",x"DD", -- 0x0208
    x"21",x"5A",x"81",x"FD",x"21",x"5A",x"81",x"32", -- 0x0210
    x"B1",x"81",x"ED",x"53",x"01",x"80",x"C3",x"65", -- 0x0218
    x"20",x"11",x"00",x"A8",x"ED",x"52",x"7D",x"01", -- 0x0220
    x"00",x"06",x"E6",x"E0",x"6F",x"7C",x"E6",x"04", -- 0x0228
    x"CA",x"39",x"22",x"CB",x"01",x"0C",x"C3",x"3B", -- 0x0230
    x"22",x"CB",x"01",x"CB",x"05",x"CB",x"14",x"10", -- 0x0238
    x"EC",x"CB",x"01",x"CB",x"01",x"CB",x"01",x"C9", -- 0x0240
    x"3A",x"CD",x"83",x"B7",x"C0",x"3A",x"04",x"80", -- 0x0248
    x"A7",x"C0",x"21",x"47",x"80",x"7E",x"4F",x"E6", -- 0x0250
    x"0F",x"FE",x"09",x"D2",x"92",x"22",x"79",x"E6", -- 0x0258
    x"F0",x"0F",x"0F",x"0F",x"0F",x"6F",x"26",x"00", -- 0x0260
    x"01",x"72",x"22",x"29",x"09",x"4E",x"23",x"66", -- 0x0268
    x"69",x"E9",x"92",x"22",x"95",x"22",x"98",x"22", -- 0x0270
    x"9B",x"22",x"A3",x"22",x"AB",x"22",x"B3",x"22", -- 0x0278
    x"BB",x"22",x"C3",x"22",x"CB",x"22",x"D3",x"22", -- 0x0280
    x"DB",x"22",x"E3",x"22",x"EB",x"22",x"F3",x"22", -- 0x0288
    x"F6",x"22",x"C3",x"6D",x"23",x"C3",x"6D",x"23", -- 0x0290
    x"C3",x"6D",x"23",x"21",x"00",x"81",x"0E",x"3C", -- 0x0298
    x"C3",x"F9",x"22",x"21",x"09",x"81",x"0E",x"1F", -- 0x02A0
    x"C3",x"F9",x"22",x"21",x"12",x"81",x"0E",x"5C", -- 0x02A8
    x"C3",x"F9",x"22",x"21",x"1B",x"81",x"0E",x"2C", -- 0x02B0
    x"C3",x"F9",x"22",x"21",x"24",x"81",x"0E",x"2F", -- 0x02B8
    x"C3",x"F9",x"22",x"C3",x"6D",x"23",x"0E",x"17", -- 0x02C0
    x"C3",x"F9",x"22",x"21",x"36",x"81",x"0E",x"22", -- 0x02C8
    x"C3",x"F9",x"22",x"21",x"3F",x"81",x"0E",x"12", -- 0x02D0
    x"C3",x"F9",x"22",x"21",x"48",x"81",x"0E",x"12", -- 0x02D8
    x"C3",x"F9",x"22",x"21",x"51",x"81",x"0E",x"12", -- 0x02E0
    x"C3",x"F9",x"22",x"21",x"5A",x"81",x"0E",x"12", -- 0x02E8
    x"C3",x"F9",x"22",x"C3",x"6D",x"23",x"C3",x"6D", -- 0x02F0
    x"23",x"3A",x"47",x"80",x"FE",x"80",x"DA",x"22", -- 0x02F8
    x"23",x"3A",x"44",x"80",x"C6",x"03",x"57",x"81", -- 0x0300
    x"5F",x"46",x"DA",x"2A",x"23",x"23",x"7E",x"BA", -- 0x0308
    x"DA",x"3F",x"23",x"BB",x"D2",x"3F",x"23",x"3A", -- 0x0310
    x"47",x"80",x"FE",x"80",x"DA",x"6D",x"23",x"C3", -- 0x0318
    x"59",x"23",x"3A",x"44",x"80",x"C6",x"0C",x"C3", -- 0x0320
    x"06",x"23",x"23",x"7E",x"BA",x"D2",x"34",x"23", -- 0x0328
    x"BB",x"D2",x"4C",x"23",x"3A",x"47",x"80",x"FE", -- 0x0330
    x"80",x"DA",x"6D",x"23",x"C3",x"59",x"23",x"10", -- 0x0338
    x"CC",x"3A",x"47",x"80",x"FE",x"80",x"DA",x"59", -- 0x0340
    x"23",x"C3",x"6D",x"23",x"10",x"DC",x"3A",x"47", -- 0x0348
    x"80",x"FE",x"80",x"DA",x"59",x"23",x"C3",x"6D", -- 0x0350
    x"23",x"3E",x"01",x"32",x"04",x"80",x"3A",x"47", -- 0x0358
    x"80",x"FE",x"80",x"D0",x"FE",x"30",x"D8",x"3E", -- 0x0360
    x"01",x"32",x"9C",x"82",x"C9",x"3A",x"04",x"80", -- 0x0368
    x"A7",x"C0",x"21",x"47",x"80",x"7E",x"C6",x"0F", -- 0x0370
    x"4F",x"E6",x"0F",x"FE",x"05",x"DA",x"B4",x"23", -- 0x0378
    x"79",x"E6",x"F0",x"0F",x"0F",x"0F",x"0F",x"6F", -- 0x0380
    x"26",x"00",x"01",x"94",x"23",x"29",x"09",x"4E", -- 0x0388
    x"23",x"66",x"69",x"E9",x"B4",x"23",x"B7",x"23", -- 0x0390
    x"BA",x"23",x"BD",x"23",x"C5",x"23",x"CD",x"23", -- 0x0398
    x"D5",x"23",x"DD",x"23",x"E5",x"23",x"ED",x"23", -- 0x03A0
    x"F5",x"23",x"FD",x"23",x"05",x"24",x"0D",x"24", -- 0x03A8
    x"15",x"24",x"15",x"24",x"C3",x"6A",x"24",x"C3", -- 0x03B0
    x"6A",x"24",x"C3",x"6A",x"24",x"21",x"00",x"81", -- 0x03B8
    x"0E",x"3C",x"C3",x"18",x"24",x"21",x"09",x"81", -- 0x03C0
    x"0E",x"1F",x"C3",x"18",x"24",x"21",x"12",x"81", -- 0x03C8
    x"0E",x"5C",x"C3",x"18",x"24",x"21",x"1B",x"81", -- 0x03D0
    x"0E",x"2C",x"C3",x"18",x"24",x"21",x"24",x"81", -- 0x03D8
    x"0E",x"2F",x"C3",x"18",x"24",x"C3",x"6A",x"24", -- 0x03E0
    x"0E",x"17",x"C3",x"18",x"24",x"21",x"36",x"81", -- 0x03E8
    x"0E",x"22",x"C3",x"18",x"24",x"21",x"3F",x"81", -- 0x03F0
    x"0E",x"12",x"C3",x"18",x"24",x"21",x"48",x"81", -- 0x03F8
    x"0E",x"12",x"C3",x"18",x"24",x"21",x"51",x"81", -- 0x0400
    x"0E",x"12",x"C3",x"18",x"24",x"21",x"5A",x"81", -- 0x0408
    x"0E",x"12",x"C3",x"18",x"24",x"C3",x"6A",x"24", -- 0x0410
    x"3A",x"2F",x"80",x"FE",x"80",x"DA",x"42",x"24", -- 0x0418
    x"3A",x"44",x"80",x"C6",x"03",x"57",x"81",x"5F", -- 0x0420
    x"46",x"DA",x"4A",x"24",x"23",x"7E",x"BA",x"DA", -- 0x0428
    x"60",x"24",x"BB",x"D2",x"60",x"24",x"3A",x"47", -- 0x0430
    x"80",x"FE",x"80",x"D8",x"3E",x"01",x"32",x"04", -- 0x0438
    x"80",x"C9",x"3A",x"44",x"80",x"C6",x"0C",x"C3", -- 0x0440
    x"25",x"24",x"23",x"7E",x"BA",x"D2",x"54",x"24", -- 0x0448
    x"BB",x"D2",x"6B",x"24",x"3A",x"47",x"80",x"FE", -- 0x0450
    x"80",x"D8",x"3E",x"01",x"32",x"04",x"80",x"C9", -- 0x0458
    x"10",x"CA",x"3A",x"47",x"80",x"FE",x"80",x"DA", -- 0x0460
    x"59",x"23",x"C9",x"10",x"DD",x"3A",x"47",x"80", -- 0x0468
    x"FE",x"80",x"DA",x"59",x"23",x"C9",x"06",x"A8", -- 0x0470
    x"08",x"A8",x"0A",x"A8",x"0C",x"A8",x"0E",x"A8", -- 0x0478
    x"10",x"A8",x"12",x"A8",x"14",x"A8",x"16",x"A8", -- 0x0480
    x"18",x"A8",x"1A",x"A8",x"5C",x"5D",x"5E",x"5F", -- 0x0488
    x"58",x"59",x"5A",x"5B",x"58",x"59",x"5A",x"5B", -- 0x0490
    x"54",x"55",x"56",x"57",x"10",x"10",x"10",x"10", -- 0x0498
    x"D0",x"D1",x"D2",x"D3",x"CC",x"CD",x"CE",x"CF", -- 0x04A0
    x"C8",x"C9",x"CA",x"CB",x"34",x"35",x"36",x"37", -- 0x04A8
    x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B", -- 0x04B0
    x"38",x"39",x"3A",x"3B",x"3C",x"3D",x"3E",x"3F", -- 0x04B8
    x"3C",x"3D",x"3E",x"3F",x"5C",x"5D",x"5E",x"5F", -- 0x04C0
    x"58",x"59",x"5A",x"5B",x"58",x"59",x"5A",x"5B", -- 0x04C8
    x"58",x"59",x"5A",x"5B",x"58",x"59",x"5A",x"5B", -- 0x04D0
    x"54",x"55",x"56",x"57",x"5C",x"5D",x"5E",x"5F", -- 0x04D8
    x"58",x"59",x"5A",x"5B",x"54",x"55",x"56",x"57", -- 0x04E0
    x"34",x"35",x"36",x"37",x"34",x"35",x"36",x"37", -- 0x04E8
    x"34",x"35",x"36",x"37",x"34",x"35",x"36",x"37", -- 0x04F0
    x"34",x"35",x"36",x"37",x"38",x"39",x"3A",x"3B", -- 0x04F8
    x"38",x"39",x"3A",x"3B",x"38",x"39",x"3A",x"3B", -- 0x0500
    x"38",x"39",x"3A",x"3B",x"38",x"39",x"3A",x"3B", -- 0x0508
    x"3C",x"3D",x"3E",x"3F",x"3C",x"3D",x"3E",x"3F", -- 0x0510
    x"3C",x"3D",x"3E",x"3F",x"3C",x"3D",x"3E",x"3F", -- 0x0518
    x"3C",x"3D",x"3E",x"3F",x"47",x"47",x"47",x"47", -- 0x0520
    x"AC",x"AD",x"AE",x"AF",x"A8",x"A9",x"AA",x"AB", -- 0x0528
    x"A0",x"A1",x"A2",x"A3",x"30",x"31",x"32",x"33", -- 0x0530
    x"A4",x"A5",x"A6",x"A7",x"50",x"51",x"52",x"53", -- 0x0538
    x"3A",x"FF",x"80",x"01",x"50",x"25",x"26",x"00", -- 0x0540
    x"87",x"6F",x"09",x"4E",x"23",x"66",x"69",x"E9", -- 0x0548
    x"66",x"25",x"77",x"25",x"88",x"25",x"99",x"25", -- 0x0550
    x"AA",x"25",x"BB",x"25",x"CC",x"25",x"DD",x"25", -- 0x0558
    x"EE",x"25",x"FF",x"25",x"10",x"26",x"21",x"9B", -- 0x0560
    x"81",x"11",x"00",x"81",x"DD",x"21",x"0C",x"80", -- 0x0568
    x"FD",x"21",x"A6",x"81",x"C3",x"21",x"26",x"21", -- 0x0570
    x"9C",x"81",x"11",x"09",x"81",x"DD",x"21",x"10", -- 0x0578
    x"80",x"FD",x"21",x"A7",x"81",x"C3",x"C7",x"26", -- 0x0580
    x"21",x"9D",x"81",x"11",x"12",x"81",x"DD",x"21", -- 0x0588
    x"14",x"80",x"FD",x"21",x"A8",x"81",x"C3",x"21", -- 0x0590
    x"26",x"21",x"9E",x"81",x"11",x"1B",x"81",x"DD", -- 0x0598
    x"21",x"18",x"80",x"FD",x"21",x"A9",x"81",x"C3", -- 0x05A0
    x"21",x"26",x"21",x"9F",x"81",x"11",x"24",x"81", -- 0x05A8
    x"DD",x"21",x"1C",x"80",x"FD",x"21",x"AA",x"81", -- 0x05B0
    x"C3",x"C7",x"26",x"C3",x"67",x"26",x"11",x"2D", -- 0x05B8
    x"81",x"DD",x"21",x"20",x"80",x"FD",x"21",x"AB", -- 0x05C0
    x"81",x"C3",x"21",x"26",x"21",x"A1",x"81",x"11", -- 0x05C8
    x"36",x"81",x"DD",x"21",x"24",x"80",x"FD",x"21", -- 0x05D0
    x"AC",x"81",x"C3",x"C7",x"26",x"21",x"A2",x"81", -- 0x05D8
    x"11",x"3F",x"81",x"DD",x"21",x"28",x"80",x"FD", -- 0x05E0
    x"21",x"AD",x"81",x"C3",x"21",x"26",x"21",x"A3", -- 0x05E8
    x"81",x"11",x"48",x"81",x"DD",x"21",x"2C",x"80", -- 0x05F0
    x"FD",x"21",x"AE",x"81",x"C3",x"C7",x"26",x"21", -- 0x05F8
    x"A4",x"81",x"11",x"51",x"81",x"DD",x"21",x"30", -- 0x0600
    x"80",x"FD",x"21",x"AF",x"81",x"C3",x"21",x"26", -- 0x0608
    x"21",x"A5",x"81",x"11",x"5A",x"81",x"DD",x"21", -- 0x0610
    x"34",x"80",x"FD",x"21",x"B0",x"81",x"C3",x"C7", -- 0x0618
    x"26",x"FD",x"7E",x"00",x"4F",x"A7",x"C2",x"5D", -- 0x0620
    x"27",x"7E",x"47",x"E6",x"0F",x"4F",x"78",x"E6", -- 0x0628
    x"10",x"C2",x"5D",x"27",x"1A",x"47",x"13",x"1A", -- 0x0630
    x"81",x"12",x"10",x"FA",x"DD",x"7E",x"00",x"81", -- 0x0638
    x"DD",x"77",x"00",x"DD",x"77",x"02",x"3A",x"47", -- 0x0640
    x"80",x"FE",x"30",x"DA",x"63",x"26",x"3A",x"47", -- 0x0648
    x"80",x"FE",x"73",x"D2",x"63",x"26",x"47",x"E6", -- 0x0650
    x"0F",x"FE",x"03",x"DA",x"74",x"26",x"FE",x"0C", -- 0x0658
    x"D2",x"A8",x"26",x"FD",x"36",x"00",x"00",x"21", -- 0x0660
    x"FF",x"80",x"34",x"7E",x"FE",x"0B",x"DA",x"40", -- 0x0668
    x"25",x"36",x"00",x"C9",x"78",x"E6",x"F0",x"08", -- 0x0670
    x"08",x"D6",x"30",x"0F",x"0F",x"0F",x"0F",x"47", -- 0x0678
    x"3A",x"FF",x"80",x"B8",x"C2",x"63",x"26",x"3A", -- 0x0680
    x"47",x"80",x"FE",x"30",x"DA",x"63",x"26",x"3A", -- 0x0688
    x"44",x"80",x"81",x"32",x"44",x"80",x"FE",x"08", -- 0x0690
    x"DA",x"A0",x"26",x"FE",x"E7",x"DA",x"63",x"26", -- 0x0698
    x"3E",x"01",x"32",x"04",x"80",x"C3",x"63",x"26", -- 0x06A0
    x"78",x"E6",x"F0",x"C6",x"10",x"08",x"08",x"D6", -- 0x06A8
    x"30",x"0F",x"0F",x"0F",x"0F",x"47",x"3A",x"FF", -- 0x06B0
    x"80",x"B8",x"C2",x"63",x"26",x"3A",x"44",x"80", -- 0x06B8
    x"81",x"32",x"44",x"80",x"C3",x"63",x"26",x"FD", -- 0x06C0
    x"7E",x"00",x"4F",x"A7",x"C2",x"6F",x"27",x"7E", -- 0x06C8
    x"47",x"E6",x"0F",x"4F",x"78",x"E6",x"10",x"C2", -- 0x06D0
    x"6F",x"27",x"1A",x"47",x"13",x"1A",x"91",x"12", -- 0x06D8
    x"10",x"FA",x"DD",x"7E",x"00",x"91",x"DD",x"77", -- 0x06E0
    x"00",x"DD",x"77",x"02",x"3A",x"47",x"80",x"FE", -- 0x06E8
    x"73",x"D2",x"01",x"27",x"47",x"E6",x"0F",x"FE", -- 0x06F0
    x"03",x"DA",x"12",x"27",x"FE",x"0C",x"D2",x"3E", -- 0x06F8
    x"27",x"FD",x"36",x"00",x"00",x"21",x"FF",x"80", -- 0x0700
    x"34",x"7E",x"FE",x"0B",x"DA",x"40",x"25",x"36", -- 0x0708
    x"00",x"C9",x"78",x"E6",x"F0",x"08",x"08",x"D6", -- 0x0710
    x"30",x"0F",x"0F",x"0F",x"0F",x"47",x"3A",x"FF", -- 0x0718
    x"80",x"B8",x"C2",x"01",x"27",x"3A",x"44",x"80", -- 0x0720
    x"91",x"32",x"44",x"80",x"FE",x"08",x"DA",x"36", -- 0x0728
    x"27",x"FE",x"E7",x"DA",x"01",x"27",x"3E",x"01", -- 0x0730
    x"32",x"04",x"80",x"C3",x"01",x"27",x"78",x"E6", -- 0x0738
    x"F0",x"C6",x"10",x"08",x"08",x"D6",x"30",x"0F", -- 0x0740
    x"0F",x"0F",x"0F",x"47",x"3A",x"FF",x"80",x"B8", -- 0x0748
    x"C2",x"01",x"27",x"3A",x"44",x"80",x"91",x"32", -- 0x0750
    x"44",x"80",x"C3",x"01",x"27",x"79",x"FE",x"01", -- 0x0758
    x"C2",x"68",x"27",x"0E",x"01",x"C3",x"34",x"26", -- 0x0760
    x"0D",x"FD",x"71",x"00",x"C3",x"67",x"26",x"79", -- 0x0768
    x"FE",x"01",x"C2",x"7A",x"27",x"0E",x"01",x"C3", -- 0x0770
    x"DA",x"26",x"0D",x"FD",x"71",x"00",x"C3",x"05", -- 0x0778
    x"27",x"3A",x"04",x"80",x"A7",x"C8",x"3A",x"50", -- 0x0780
    x"81",x"CB",x"47",x"28",x"05",x"3E",x"01",x"32", -- 0x0788
    x"18",x"81",x"3A",x"20",x"81",x"A7",x"28",x"03", -- 0x0790
    x"32",x"21",x"81",x"CD",x"57",x"36",x"CD",x"3C", -- 0x0798
    x"38",x"3A",x"47",x"82",x"3C",x"32",x"47",x"82", -- 0x07A0
    x"D6",x"10",x"C0",x"32",x"47",x"82",x"3E",x"07", -- 0x07A8
    x"32",x"46",x"80",x"21",x"44",x"80",x"3A",x"B2", -- 0x07B0
    x"81",x"3C",x"32",x"B2",x"81",x"4F",x"3A",x"9C", -- 0x07B8
    x"82",x"A7",x"C2",x"06",x"28",x"79",x"FE",x"06", -- 0x07C0
    x"20",x"44",x"CD",x"17",x"08",x"AF",x"32",x"B2", -- 0x07C8
    x"81",x"32",x"04",x"80",x"32",x"47",x"82",x"32", -- 0x07D0
    x"69",x"82",x"32",x"9C",x"82",x"21",x"48",x"82", -- 0x07D8
    x"11",x"49",x"82",x"01",x"0B",x"00",x"77",x"ED", -- 0x07E0
    x"B0",x"3C",x"32",x"CE",x"83",x"3A",x"D6",x"83", -- 0x07E8
    x"3D",x"20",x"12",x"3A",x"FE",x"83",x"A7",x"20", -- 0x07F0
    x"0C",x"32",x"D6",x"83",x"32",x"99",x"82",x"32", -- 0x07F8
    x"9A",x"82",x"32",x"5B",x"82",x"C9",x"79",x"FE", -- 0x0800
    x"05",x"20",x"03",x"C3",x"CA",x"27",x"3A",x"9C", -- 0x0808
    x"82",x"A7",x"C2",x"4D",x"28",x"23",x"3A",x"B2", -- 0x0810
    x"81",x"3D",x"28",x"0B",x"3D",x"28",x"15",x"3D", -- 0x0818
    x"28",x"15",x"3D",x"28",x"15",x"18",x"16",x"36", -- 0x0820
    x"39",x"AF",x"67",x"6F",x"22",x"82",x"83",x"DF", -- 0x0828
    x"3E",x"03",x"DF",x"C9",x"36",x"39",x"C9",x"36", -- 0x0830
    x"3A",x"C9",x"36",x"3B",x"C9",x"36",x"3C",x"AF", -- 0x0838
    x"32",x"AE",x"83",x"CD",x"DF",x"38",x"21",x"D8", -- 0x0840
    x"00",x"22",x"82",x"83",x"C9",x"23",x"3A",x"B2", -- 0x0848
    x"81",x"3D",x"28",x"08",x"3D",x"28",x"12",x"3D", -- 0x0850
    x"28",x"12",x"18",x"13",x"36",x"22",x"AF",x"67", -- 0x0858
    x"6F",x"22",x"82",x"83",x"DF",x"3E",x"02",x"DF", -- 0x0860
    x"C9",x"36",x"23",x"C9",x"36",x"24",x"C9",x"36", -- 0x0868
    x"3C",x"AF",x"32",x"AE",x"83",x"32",x"10",x"81", -- 0x0870
    x"32",x"07",x"81",x"32",x"1A",x"81",x"32",x"19", -- 0x0878
    x"81",x"CD",x"DF",x"38",x"21",x"D8",x"00",x"22", -- 0x0880
    x"82",x"83",x"C9",x"3A",x"4F",x"81",x"A7",x"C0", -- 0x0888
    x"3A",x"5B",x"81",x"A7",x"C0",x"3A",x"B4",x"81", -- 0x0890
    x"A7",x"C2",x"BB",x"28",x"67",x"3A",x"B3",x"81", -- 0x0898
    x"6F",x"11",x"CA",x"28",x"29",x"19",x"4E",x"23", -- 0x08A0
    x"66",x"69",x"EB",x"21",x"B3",x"81",x"34",x"7E", -- 0x08A8
    x"23",x"36",x"15",x"D6",x"0A",x"C2",x"C0",x"28", -- 0x08B0
    x"2B",x"77",x"C9",x"21",x"B4",x"81",x"35",x"C9", -- 0x08B8
    x"EB",x"11",x"9B",x"81",x"01",x"0B",x"00",x"ED", -- 0x08C0
    x"B0",x"C9",x"F4",x"28",x"FF",x"28",x"0A",x"29", -- 0x08C8
    x"15",x"29",x"20",x"29",x"2B",x"29",x"36",x"29", -- 0x08D0
    x"41",x"29",x"4C",x"29",x"57",x"29",x"62",x"29", -- 0x08D8
    x"6D",x"29",x"78",x"29",x"83",x"29",x"8E",x"29", -- 0x08E0
    x"99",x"29",x"A4",x"29",x"AF",x"29",x"BA",x"29", -- 0x08E8
    x"C5",x"29",x"D0",x"29",x"13",x"12",x"11",x"16", -- 0x08F0
    x"12",x"00",x"12",x"13",x"14",x"15",x"16",x"12", -- 0x08F8
    x"13",x"12",x"15",x"01",x"00",x"13",x"02",x"12", -- 0x0900
    x"13",x"12",x"12",x"12",x"13",x"14",x"12",x"00", -- 0x0908
    x"12",x"01",x"13",x"12",x"13",x"12",x"01",x"12", -- 0x0910
    x"13",x"13",x"00",x"12",x"02",x"12",x"01",x"14", -- 0x0918
    x"13",x"12",x"01",x"12",x"12",x"00",x"12",x"01", -- 0x0920
    x"01",x"12",x"13",x"13",x"01",x"12",x"13",x"13", -- 0x0928
    x"00",x"01",x"02",x"12",x"13",x"12",x"12",x"12", -- 0x0930
    x"13",x"12",x"12",x"00",x"12",x"01",x"13",x"12", -- 0x0938
    x"13",x"13",x"13",x"12",x"13",x"01",x"00",x"13", -- 0x0940
    x"02",x"12",x"01",x"12",x"12",x"12",x"13",x"12", -- 0x0948
    x"12",x"00",x"12",x"01",x"01",x"12",x"13",x"13", -- 0x0950
    x"01",x"12",x"01",x"13",x"00",x"01",x"02",x"12", -- 0x0958
    x"13",x"13",x"12",x"12",x"01",x"12",x"12",x"00", -- 0x0960
    x"01",x"01",x"13",x"12",x"12",x"01",x"13",x"01", -- 0x0968
    x"13",x"01",x"00",x"12",x"01",x"12",x"01",x"01", -- 0x0970
    x"12",x"12",x"01",x"12",x"12",x"00",x"01",x"02", -- 0x0978
    x"13",x"12",x"01",x"01",x"12",x"01",x"12",x"01", -- 0x0980
    x"00",x"01",x"03",x"12",x"01",x"12",x"12",x"12", -- 0x0988
    x"01",x"12",x"12",x"00",x"01",x"02",x"13",x"12", -- 0x0990
    x"12",x"01",x"01",x"12",x"01",x"12",x"00",x"01", -- 0x0998
    x"01",x"12",x"01",x"01",x"01",x"01",x"12",x"01", -- 0x09A0
    x"12",x"00",x"01",x"01",x"12",x"01",x"01",x"12", -- 0x09A8
    x"01",x"13",x"12",x"01",x"00",x"12",x"02",x"01", -- 0x09B0
    x"12",x"12",x"01",x"12",x"14",x"01",x"12",x"00", -- 0x09B8
    x"01",x"03",x"12",x"13",x"01",x"12",x"01",x"13", -- 0x09C0
    x"12",x"13",x"00",x"12",x"02",x"13",x"12",x"12", -- 0x09C8
    x"13",x"12",x"12",x"13",x"12",x"00",x"13",x"01", -- 0x09D0
    x"14",x"13",x"14",x"21",x"43",x"A8",x"0E",x"05", -- 0x09D8
    x"11",x"7F",x"2A",x"06",x"04",x"1A",x"77",x"13", -- 0x09E0
    x"C5",x"01",x"20",x"00",x"09",x"C1",x"10",x"F5", -- 0x09E8
    x"11",x"40",x"00",x"19",x"0D",x"C2",x"E0",x"29", -- 0x09F0
    x"21",x"A4",x"A8",x"0E",x"04",x"11",x"83",x"2A", -- 0x09F8
    x"06",x"04",x"1A",x"77",x"13",x"C5",x"01",x"20", -- 0x0A00
    x"00",x"09",x"C1",x"10",x"F5",x"11",x"40",x"00", -- 0x0A08
    x"19",x"0D",x"C2",x"FD",x"29",x"21",x"A5",x"A8", -- 0x0A10
    x"0E",x"04",x"11",x"87",x"2A",x"06",x"04",x"1A", -- 0x0A18
    x"77",x"13",x"C5",x"01",x"20",x"00",x"09",x"C1", -- 0x0A20
    x"10",x"F5",x"11",x"40",x"00",x"19",x"0D",x"C2", -- 0x0A28
    x"1A",x"2A",x"21",x"C3",x"A8",x"06",x"04",x"36", -- 0x0A30
    x"47",x"11",x"20",x"00",x"19",x"36",x"47",x"11", -- 0x0A38
    x"A0",x"00",x"19",x"10",x"F2",x"21",x"44",x"A8", -- 0x0A40
    x"36",x"41",x"23",x"36",x"42",x"01",x"5F",x"03", -- 0x0A48
    x"09",x"36",x"45",x"23",x"36",x"46",x"21",x"5C", -- 0x0A50
    x"A8",x"CD",x"6B",x"2A",x"21",x"07",x"80",x"3E", -- 0x0A58
    x"01",x"77",x"2C",x"2C",x"77",x"2C",x"2C",x"77", -- 0x0A60
    x"C3",x"8B",x"2A",x"06",x"0E",x"36",x"48",x"23", -- 0x0A68
    x"36",x"49",x"11",x"1F",x"00",x"19",x"36",x"4A", -- 0x0A70
    x"23",x"36",x"4B",x"19",x"10",x"EF",x"C9",x"40", -- 0x0A78
    x"43",x"43",x"44",x"45",x"47",x"47",x"41",x"46", -- 0x0A80
    x"43",x"43",x"42",x"3E",x"05",x"32",x"25",x"80", -- 0x0A88
    x"32",x"27",x"80",x"3E",x"04",x"32",x"2D",x"80", -- 0x0A90
    x"32",x"2F",x"80",x"3E",x"07",x"32",x"35",x"80", -- 0x0A98
    x"32",x"37",x"80",x"3E",x"06",x"32",x"21",x"80", -- 0x0AA0
    x"32",x"23",x"80",x"32",x"39",x"80",x"32",x"3B", -- 0x0AA8
    x"80",x"3E",x"05",x"06",x"0A",x"21",x"0D",x"80", -- 0x0AB0
    x"77",x"23",x"23",x"10",x"FB",x"32",x"29",x"80", -- 0x0AB8
    x"32",x"2B",x"80",x"32",x"31",x"80",x"32",x"33", -- 0x0AC0
    x"80",x"3E",x"02",x"32",x"0D",x"80",x"32",x"0F", -- 0x0AC8
    x"80",x"32",x"15",x"80",x"32",x"17",x"80",x"32", -- 0x0AD0
    x"19",x"80",x"32",x"1B",x"80",x"C9",x"3A",x"FE", -- 0x0AD8
    x"83",x"B7",x"28",x"34",x"CD",x"44",x"39",x"CD", -- 0x0AE0
    x"A6",x"39",x"CD",x"73",x"38",x"CD",x"2F",x"37", -- 0x0AE8
    x"CD",x"8F",x"39",x"3A",x"40",x"83",x"A7",x"C4", -- 0x0AF0
    x"28",x"2B",x"CD",x"74",x"34",x"3A",x"B7",x"83", -- 0x0AF8
    x"CB",x"47",x"CA",x"36",x"2B",x"3A",x"22",x"81", -- 0x0B00
    x"3C",x"32",x"22",x"81",x"A7",x"CC",x"83",x"34", -- 0x0B08
    x"3A",x"22",x"81",x"FE",x"70",x"CC",x"57",x"36", -- 0x0B10
    x"3A",x"47",x"80",x"FE",x"31",x"DA",x"88",x"2D", -- 0x0B18
    x"3A",x"FE",x"83",x"B7",x"C8",x"C3",x"54",x"2B", -- 0x0B20
    x"3D",x"32",x"40",x"83",x"FE",x"01",x"C0",x"CD", -- 0x0B28
    x"23",x"37",x"CD",x"67",x"38",x"C9",x"3A",x"22", -- 0x0B30
    x"81",x"3C",x"32",x"22",x"81",x"A7",x"CC",x"1F", -- 0x0B38
    x"35",x"3A",x"22",x"81",x"FE",x"50",x"CC",x"BB", -- 0x0B40
    x"35",x"3A",x"22",x"81",x"FE",x"B0",x"CC",x"57", -- 0x0B48
    x"36",x"C3",x"18",x"2B",x"3A",x"6C",x"82",x"A7", -- 0x0B50
    x"C0",x"3A",x"68",x"82",x"A7",x"28",x"08",x"3D", -- 0x0B58
    x"32",x"68",x"82",x"CD",x"74",x"34",x"C9",x"3A", -- 0x0B60
    x"04",x"80",x"A7",x"C0",x"21",x"44",x"80",x"11", -- 0x0B68
    x"47",x"80",x"3A",x"04",x"E0",x"CB",x"5F",x"28", -- 0x0B70
    x"07",x"3A",x"FD",x"83",x"3D",x"C2",x"FD",x"2B", -- 0x0B78
    x"3A",x"00",x"E0",x"4F",x"3A",x"48",x"82",x"A7", -- 0x0B80
    x"C2",x"43",x"2C",x"3A",x"04",x"E0",x"CB",x"5F", -- 0x0B88
    x"28",x"07",x"3A",x"FD",x"83",x"3D",x"C2",x"04", -- 0x0B90
    x"2C",x"3A",x"04",x"E0",x"CB",x"77",x"CA",x"14", -- 0x0B98
    x"2C",x"AF",x"32",x"4C",x"82",x"32",x"50",x"82", -- 0x0BA0
    x"3A",x"49",x"82",x"A7",x"C2",x"96",x"2C",x"3A", -- 0x0BA8
    x"4A",x"82",x"47",x"3A",x"4B",x"82",x"80",x"20", -- 0x0BB0
    x"1D",x"3A",x"04",x"E0",x"CB",x"5F",x"28",x"07", -- 0x0BB8
    x"3A",x"FD",x"83",x"3D",x"C2",x"0C",x"2C",x"3A", -- 0x0BC0
    x"04",x"E0",x"CB",x"67",x"CA",x"6D",x"2C",x"AF", -- 0x0BC8
    x"32",x"4D",x"82",x"32",x"51",x"82",x"3A",x"4A", -- 0x0BD0
    x"82",x"A7",x"C2",x"FF",x"2C",x"CB",x"61",x"CA", -- 0x0BD8
    x"CA",x"2C",x"AF",x"32",x"4E",x"82",x"32",x"52", -- 0x0BE0
    x"82",x"3A",x"4B",x"82",x"A7",x"C2",x"5E",x"2D", -- 0x0BE8
    x"CB",x"69",x"CA",x"29",x"2D",x"AF",x"32",x"4F", -- 0x0BF0
    x"82",x"32",x"53",x"82",x"C9",x"3A",x"02",x"E0", -- 0x0BF8
    x"4F",x"C3",x"84",x"2B",x"3A",x"04",x"E0",x"CB", -- 0x0C00
    x"47",x"C3",x"9E",x"2B",x"3A",x"00",x"E0",x"CB", -- 0x0C08
    x"47",x"C3",x"CC",x"2B",x"3A",x"47",x"80",x"FE", -- 0x0C10
    x"F0",x"D0",x"3A",x"50",x"82",x"A7",x"20",x"10", -- 0x0C18
    x"3E",x"04",x"DF",x"23",x"7E",x"2B",x"FE",x"DE", -- 0x0C20
    x"CA",x"3D",x"2C",x"3E",x"DE",x"32",x"45",x"80", -- 0x0C28
    x"3A",x"50",x"82",x"3C",x"32",x"50",x"82",x"B7", -- 0x0C30
    x"C8",x"AF",x"32",x"50",x"82",x"3A",x"56",x"82", -- 0x0C38
    x"32",x"50",x"82",x"3A",x"4C",x"82",x"A7",x"C0", -- 0x0C40
    x"3C",x"32",x"48",x"82",x"3A",x"50",x"82",x"3D", -- 0x0C48
    x"32",x"50",x"82",x"C2",x"61",x"2C",x"32",x"48", -- 0x0C50
    x"82",x"3C",x"32",x"4C",x"82",x"23",x"36",x"DE", -- 0x0C58
    x"C9",x"EB",x"3A",x"54",x"82",x"86",x"77",x"EB", -- 0x0C60
    x"23",x"3E",x"DC",x"77",x"C9",x"3A",x"51",x"82", -- 0x0C68
    x"A7",x"20",x"10",x"3E",x"04",x"DF",x"23",x"7E", -- 0x0C70
    x"2B",x"FE",x"1E",x"CA",x"90",x"2C",x"3E",x"1E", -- 0x0C78
    x"32",x"45",x"80",x"3A",x"51",x"82",x"3C",x"32", -- 0x0C80
    x"51",x"82",x"B7",x"C8",x"AF",x"32",x"51",x"82", -- 0x0C88
    x"3A",x"57",x"82",x"32",x"51",x"82",x"CD",x"74", -- 0x0C90
    x"34",x"3A",x"4D",x"82",x"A7",x"C0",x"3C",x"32", -- 0x0C98
    x"49",x"82",x"3A",x"51",x"82",x"3D",x"32",x"51", -- 0x0CA0
    x"82",x"C2",x"BC",x"2C",x"32",x"49",x"82",x"3C", -- 0x0CA8
    x"32",x"4D",x"82",x"23",x"36",x"1E",x"D5",x"CD", -- 0x0CB0
    x"5F",x"30",x"D1",x"C9",x"EB",x"3A",x"54",x"82", -- 0x0CB8
    x"47",x"7E",x"90",x"77",x"EB",x"23",x"3E",x"1C", -- 0x0CC0
    x"77",x"C9",x"3A",x"47",x"80",x"FE",x"30",x"D8", -- 0x0CC8
    x"3A",x"44",x"80",x"FE",x"E0",x"D0",x"3A",x"52", -- 0x0CD0
    x"82",x"A7",x"20",x"10",x"3E",x"04",x"DF",x"23", -- 0x0CD8
    x"7E",x"2B",x"FE",x"A1",x"CA",x"F9",x"2C",x"3E", -- 0x0CE0
    x"A1",x"32",x"45",x"80",x"3A",x"52",x"82",x"3C", -- 0x0CE8
    x"32",x"52",x"82",x"B7",x"C8",x"AF",x"32",x"52", -- 0x0CF0
    x"82",x"3A",x"58",x"82",x"32",x"52",x"82",x"3A", -- 0x0CF8
    x"4E",x"82",x"A7",x"C0",x"3C",x"32",x"4A",x"82", -- 0x0D00
    x"3A",x"52",x"82",x"3D",x"32",x"52",x"82",x"C2", -- 0x0D08
    x"1D",x"2D",x"32",x"4A",x"82",x"3C",x"32",x"4E", -- 0x0D10
    x"82",x"23",x"36",x"A1",x"C9",x"3A",x"55",x"82", -- 0x0D18
    x"47",x"7E",x"80",x"77",x"23",x"3E",x"9F",x"77", -- 0x0D20
    x"C9",x"3A",x"47",x"80",x"FE",x"30",x"D8",x"3A", -- 0x0D28
    x"44",x"80",x"FE",x"20",x"D8",x"3A",x"53",x"82", -- 0x0D30
    x"A7",x"20",x"10",x"3E",x"04",x"DF",x"23",x"7E", -- 0x0D38
    x"2B",x"FE",x"21",x"CA",x"58",x"2D",x"3E",x"21", -- 0x0D40
    x"32",x"45",x"80",x"3A",x"53",x"82",x"3C",x"32", -- 0x0D48
    x"53",x"82",x"B7",x"C8",x"AF",x"32",x"53",x"82", -- 0x0D50
    x"3A",x"59",x"82",x"32",x"53",x"82",x"3A",x"4F", -- 0x0D58
    x"82",x"A7",x"C0",x"3C",x"32",x"4B",x"82",x"3A", -- 0x0D60
    x"53",x"82",x"3D",x"32",x"53",x"82",x"C2",x"7C", -- 0x0D68
    x"2D",x"32",x"4B",x"82",x"3C",x"32",x"4F",x"82", -- 0x0D70
    x"23",x"36",x"21",x"C9",x"3A",x"55",x"82",x"47", -- 0x0D78
    x"7E",x"90",x"77",x"23",x"3E",x"1F",x"77",x"C9", -- 0x0D80
    x"3A",x"44",x"80",x"FE",x"15",x"DA",x"00",x"2E", -- 0x0D88
    x"FE",x"1C",x"CA",x"10",x"2E",x"DA",x"10",x"2E", -- 0x0D90
    x"FE",x"2E",x"DA",x"00",x"2E",x"FE",x"35",x"CA", -- 0x0D98
    x"00",x"2E",x"DA",x"00",x"2E",x"FE",x"45",x"DA", -- 0x0DA0
    x"00",x"2E",x"FE",x"4C",x"CA",x"61",x"2E",x"DA", -- 0x0DA8
    x"61",x"2E",x"FE",x"5E",x"DA",x"00",x"2E",x"FE", -- 0x0DB0
    x"65",x"CA",x"00",x"2E",x"DA",x"00",x"2E",x"FE", -- 0x0DB8
    x"75",x"DA",x"00",x"2E",x"FE",x"7C",x"CA",x"B2", -- 0x0DC0
    x"2E",x"DA",x"B2",x"2E",x"FE",x"8E",x"DA",x"00", -- 0x0DC8
    x"2E",x"FE",x"95",x"CA",x"00",x"2E",x"DA",x"00", -- 0x0DD0
    x"2E",x"FE",x"A5",x"DA",x"00",x"2E",x"FE",x"AC", -- 0x0DD8
    x"CA",x"03",x"2F",x"DA",x"03",x"2F",x"FE",x"BE", -- 0x0DE0
    x"DA",x"00",x"2E",x"FE",x"C5",x"CA",x"00",x"2E", -- 0x0DE8
    x"DA",x"00",x"2E",x"FE",x"D5",x"DA",x"00",x"2E", -- 0x0DF0
    x"FE",x"DC",x"CA",x"54",x"2F",x"DA",x"54",x"2F", -- 0x0DF8
    x"3A",x"47",x"80",x"FE",x"2A",x"D2",x"54",x"2B", -- 0x0E00
    x"3E",x"01",x"32",x"04",x"80",x"C3",x"54",x"2B", -- 0x0E08
    x"3A",x"FD",x"83",x"3D",x"20",x"3C",x"3A",x"5E", -- 0x0E10
    x"82",x"A7",x"C0",x"3A",x"47",x"80",x"FE",x"2A", -- 0x0E18
    x"D2",x"54",x"2B",x"06",x"18",x"3A",x"21",x"81", -- 0x0E20
    x"D6",x"01",x"CC",x"FC",x"36",x"21",x"64",x"AB", -- 0x0E28
    x"CD",x"A5",x"2F",x"3A",x"34",x"81",x"A7",x"28", -- 0x0E30
    x"09",x"06",x"18",x"CD",x"54",x"38",x"AF",x"32", -- 0x0E38
    x"34",x"81",x"3A",x"FD",x"83",x"3D",x"20",x"0F", -- 0x0E40
    x"3E",x"01",x"32",x"5E",x"82",x"21",x"5C",x"82", -- 0x0E48
    x"34",x"C9",x"3A",x"63",x"82",x"18",x"C2",x"3E", -- 0x0E50
    x"01",x"32",x"63",x"82",x"21",x"5D",x"82",x"34", -- 0x0E58
    x"C9",x"3A",x"FD",x"83",x"3D",x"20",x"3C",x"3A", -- 0x0E60
    x"5F",x"82",x"A7",x"C0",x"3A",x"47",x"80",x"FE", -- 0x0E68
    x"2A",x"D2",x"54",x"2B",x"06",x"48",x"3A",x"21", -- 0x0E70
    x"81",x"D6",x"02",x"CC",x"FC",x"36",x"21",x"A4", -- 0x0E78
    x"AA",x"CD",x"A5",x"2F",x"3A",x"34",x"81",x"A7", -- 0x0E80
    x"28",x"09",x"06",x"48",x"CD",x"54",x"38",x"AF", -- 0x0E88
    x"32",x"34",x"81",x"3A",x"FD",x"83",x"3D",x"20", -- 0x0E90
    x"0F",x"3E",x"01",x"32",x"5F",x"82",x"21",x"5C", -- 0x0E98
    x"82",x"34",x"C9",x"3A",x"64",x"82",x"18",x"C2", -- 0x0EA0
    x"3E",x"01",x"32",x"64",x"82",x"21",x"5D",x"82", -- 0x0EA8
    x"34",x"C9",x"3A",x"FD",x"83",x"3D",x"20",x"3C", -- 0x0EB0
    x"3A",x"60",x"82",x"A7",x"C0",x"3A",x"47",x"80", -- 0x0EB8
    x"FE",x"2A",x"D2",x"54",x"2B",x"06",x"78",x"3A", -- 0x0EC0
    x"21",x"81",x"D6",x"03",x"CC",x"FC",x"36",x"21", -- 0x0EC8
    x"E4",x"A9",x"CD",x"A5",x"2F",x"3A",x"34",x"81", -- 0x0ED0
    x"A7",x"28",x"09",x"06",x"78",x"CD",x"54",x"38", -- 0x0ED8
    x"AF",x"32",x"34",x"81",x"3A",x"FD",x"83",x"3D", -- 0x0EE0
    x"20",x"0F",x"3E",x"01",x"32",x"60",x"82",x"21", -- 0x0EE8
    x"5C",x"82",x"34",x"C9",x"3A",x"65",x"82",x"18", -- 0x0EF0
    x"C2",x"3E",x"01",x"32",x"65",x"82",x"21",x"5D", -- 0x0EF8
    x"82",x"34",x"C9",x"3A",x"FD",x"83",x"3D",x"20", -- 0x0F00
    x"3C",x"3A",x"61",x"82",x"A7",x"C0",x"3A",x"47", -- 0x0F08
    x"80",x"FE",x"2A",x"D2",x"54",x"2B",x"06",x"A8", -- 0x0F10
    x"3A",x"21",x"81",x"D6",x"04",x"CC",x"FC",x"36", -- 0x0F18
    x"21",x"24",x"A9",x"CD",x"A5",x"2F",x"3A",x"34", -- 0x0F20
    x"81",x"A7",x"28",x"09",x"06",x"A8",x"CD",x"54", -- 0x0F28
    x"38",x"AF",x"32",x"34",x"81",x"3A",x"FD",x"83", -- 0x0F30
    x"3D",x"20",x"0F",x"3E",x"01",x"32",x"61",x"82", -- 0x0F38
    x"21",x"5C",x"82",x"34",x"C9",x"3A",x"66",x"82", -- 0x0F40
    x"18",x"C2",x"3E",x"01",x"32",x"66",x"82",x"21", -- 0x0F48
    x"5D",x"82",x"34",x"C9",x"3A",x"FD",x"83",x"3D", -- 0x0F50
    x"20",x"3C",x"3A",x"62",x"82",x"A7",x"C0",x"3A", -- 0x0F58
    x"47",x"80",x"FE",x"2A",x"D2",x"54",x"2B",x"06", -- 0x0F60
    x"D8",x"3A",x"21",x"81",x"D6",x"05",x"CC",x"FC", -- 0x0F68
    x"36",x"21",x"64",x"A8",x"CD",x"A5",x"2F",x"3A", -- 0x0F70
    x"34",x"81",x"A7",x"28",x"09",x"06",x"D8",x"CD", -- 0x0F78
    x"54",x"38",x"AF",x"32",x"34",x"81",x"3A",x"FD", -- 0x0F80
    x"83",x"3D",x"20",x"0F",x"3E",x"01",x"32",x"62", -- 0x0F88
    x"82",x"21",x"5C",x"82",x"34",x"C9",x"3A",x"67", -- 0x0F90
    x"82",x"18",x"C2",x"3E",x"01",x"32",x"67",x"82", -- 0x0F98
    x"21",x"5D",x"82",x"34",x"C9",x"3A",x"34",x"81", -- 0x0FA0
    x"A7",x"28",x"09",x"11",x"20",x"00",x"CD",x"03", -- 0x0FA8
    x"09",x"CD",x"45",x"38",x"36",x"6C",x"23",x"36", -- 0x0FB0
    x"6D",x"01",x"1F",x"00",x"09",x"36",x"6E",x"23", -- 0x0FB8
    x"36",x"6F",x"E5",x"D5",x"11",x"05",x"00",x"CD", -- 0x0FC0
    x"03",x"09",x"CD",x"E8",x"08",x"3A",x"FE",x"83", -- 0x0FC8
    x"B7",x"28",x"4A",x"AF",x"67",x"6F",x"22",x"82", -- 0x0FD0
    x"83",x"DF",x"3E",x"F0",x"DF",x"3A",x"FD",x"83", -- 0x0FD8
    x"21",x"5C",x"82",x"3D",x"28",x"01",x"2C",x"7E", -- 0x0FE0
    x"FE",x"04",x"28",x"1E",x"3E",x"08",x"DF",x"3E", -- 0x0FE8
    x"0E",x"DF",x"21",x"81",x"83",x"35",x"20",x"02", -- 0x0FF0
    x"36",x"14",x"7E",x"21",x"5D",x"0F",x"87",x"85"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
