-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity SCRAMBLE_PGM_01 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of SCRAMBLE_PGM_01 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"3A",x"00",x"40",x"FE",x"55",x"CA",x"01",x"40", -- 0x0000
    x"3A",x"00",x"88",x"31",x"00",x"88",x"C3",x"B1", -- 0x0008
    x"02",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0010
    x"4F",x"3A",x"FE",x"83",x"B7",x"C8",x"E5",x"21", -- 0x0018
    x"00",x"83",x"34",x"7E",x"6F",x"71",x"E1",x"C9", -- 0x0020
    x"1A",x"77",x"7D",x"D6",x"20",x"6F",x"30",x"01", -- 0x0028
    x"25",x"13",x"10",x"F4",x"C9",x"FF",x"FF",x"FF", -- 0x0030
    x"11",x"10",x"20",x"21",x"00",x"A8",x"06",x"20", -- 0x0038
    x"73",x"23",x"10",x"FC",x"0E",x"15",x"10",x"FE", -- 0x0040
    x"0D",x"20",x"FB",x"15",x"20",x"F0",x"C9",x"FF", -- 0x0048
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0050
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"E5", -- 0x0060
    x"D5",x"C5",x"DD",x"E5",x"FD",x"E5",x"3A",x"00", -- 0x0068
    x"88",x"AF",x"32",x"08",x"B8",x"CD",x"00",x"3E", -- 0x0070
    x"21",x"07",x"80",x"11",x"07",x"B0",x"7E",x"12", -- 0x0078
    x"2C",x"1C",x"06",x"1C",x"7E",x"0F",x"0F",x"0F", -- 0x0080
    x"0F",x"12",x"2C",x"1C",x"7E",x"12",x"2C",x"1C", -- 0x0088
    x"10",x"F2",x"0E",x"08",x"3A",x"2F",x"84",x"B7", -- 0x0090
    x"28",x"05",x"0E",x"06",x"1E",x"48",x"6B",x"7E", -- 0x0098
    x"0F",x"0F",x"0F",x"0F",x"12",x"2C",x"1C",x"06", -- 0x00A0
    x"03",x"7E",x"12",x"2C",x"1C",x"10",x"FA",x"0D", -- 0x00A8
    x"20",x"ED",x"21",x"7F",x"83",x"7E",x"B7",x"28", -- 0x00B0
    x"07",x"35",x"20",x"04",x"AF",x"32",x"1C",x"B8", -- 0x00B8
    x"21",x"7E",x"83",x"7E",x"B7",x"28",x"07",x"35", -- 0x00C0
    x"20",x"04",x"AF",x"32",x"18",x"B8",x"3A",x"04", -- 0x00C8
    x"E0",x"E6",x"08",x"CA",x"FC",x"00",x"3A",x"FE", -- 0x00D0
    x"83",x"A7",x"CA",x"FC",x"00",x"3A",x"FD",x"83", -- 0x00D8
    x"A7",x"28",x"19",x"3D",x"28",x"16",x"0E",x"02", -- 0x00E0
    x"21",x"43",x"80",x"11",x"43",x"B0",x"7E",x"81", -- 0x00E8
    x"12",x"0E",x"02",x"21",x"47",x"80",x"11",x"47", -- 0x00F0
    x"B0",x"7E",x"81",x"12",x"3A",x"FE",x"83",x"B7", -- 0x00F8
    x"CA",x"22",x"01",x"CD",x"BF",x"07",x"3A",x"EA", -- 0x0100
    x"83",x"B7",x"CA",x"53",x"02",x"2A",x"D2",x"83", -- 0x0108
    x"7C",x"B5",x"CA",x"7F",x"01",x"2B",x"22",x"D2", -- 0x0110
    x"83",x"CD",x"40",x"25",x"CD",x"8B",x"28",x"C3", -- 0x0118
    x"53",x"02",x"3A",x"86",x"83",x"A7",x"CA",x"30", -- 0x0120
    x"01",x"3D",x"32",x"86",x"83",x"C3",x"53",x"02", -- 0x0128
    x"3A",x"D6",x"83",x"FE",x"02",x"D2",x"66",x"01", -- 0x0130
    x"B7",x"CC",x"D4",x"0D",x"CD",x"CA",x"33",x"AF", -- 0x0138
    x"32",x"CD",x"83",x"32",x"CF",x"83",x"32",x"B5", -- 0x0140
    x"83",x"67",x"6F",x"22",x"93",x"82",x"21",x"5C", -- 0x0148
    x"82",x"11",x"5D",x"82",x"01",x"0B",x"00",x"70", -- 0x0150
    x"ED",x"B0",x"21",x"AF",x"83",x"36",x"80",x"2C", -- 0x0158
    x"77",x"2C",x"77",x"C3",x"53",x"02",x"21",x"D8", -- 0x0160
    x"83",x"7E",x"B7",x"CA",x"53",x"02",x"35",x"C2", -- 0x0168
    x"53",x"02",x"2D",x"7E",x"B7",x"C2",x"53",x"02", -- 0x0170
    x"21",x"D6",x"83",x"35",x"C3",x"53",x"02",x"2A", -- 0x0178
    x"82",x"83",x"7C",x"B5",x"28",x"12",x"2B",x"22", -- 0x0180
    x"82",x"83",x"7C",x"B5",x"20",x"0A",x"3E",x"0F", -- 0x0188
    x"DF",x"3E",x"B0",x"DF",x"AF",x"32",x"71",x"83", -- 0x0190
    x"3A",x"FD",x"83",x"3D",x"C2",x"82",x"02",x"3A", -- 0x0198
    x"5C",x"82",x"FE",x"05",x"CA",x"6C",x"02",x"3A", -- 0x01A0
    x"98",x"82",x"A7",x"28",x"07",x"3D",x"32",x"98", -- 0x01A8
    x"82",x"C3",x"F0",x"01",x"3A",x"97",x"82",x"A7", -- 0x01B0
    x"C2",x"65",x"02",x"2A",x"9D",x"82",x"7C",x"B5", -- 0x01B8
    x"20",x"2E",x"CD",x"93",x"08",x"CD",x"DE",x"2A", -- 0x01C0
    x"3A",x"B5",x"83",x"B7",x"20",x"22",x"3C",x"32", -- 0x01C8
    x"B5",x"83",x"3E",x"FF",x"32",x"84",x"83",x"3A", -- 0x01D0
    x"80",x"83",x"B7",x"28",x"13",x"AF",x"32",x"80", -- 0x01D8
    x"83",x"21",x"40",x"00",x"22",x"82",x"83",x"11", -- 0x01E0
    x"11",x"10",x"21",x"51",x"AA",x"06",x"07",x"EF", -- 0x01E8
    x"3A",x"84",x"83",x"B7",x"28",x"0A",x"3D",x"32", -- 0x01F0
    x"84",x"83",x"21",x"50",x"A8",x"CC",x"6B",x"2A", -- 0x01F8
    x"CD",x"8E",x"30",x"CD",x"8B",x"28",x"3A",x"07", -- 0x0200
    x"81",x"A7",x"28",x"07",x"3A",x"09",x"81",x"3D", -- 0x0208
    x"32",x"09",x"81",x"3A",x"08",x"81",x"A7",x"28", -- 0x0210
    x"07",x"3A",x"24",x"81",x"3D",x"32",x"24",x"81", -- 0x0218
    x"CD",x"48",x"22",x"3A",x"07",x"81",x"A7",x"28", -- 0x0220
    x"07",x"3A",x"09",x"81",x"3C",x"32",x"09",x"81", -- 0x0228
    x"3A",x"08",x"81",x"A7",x"28",x"07",x"3A",x"24", -- 0x0230
    x"81",x"3C",x"32",x"24",x"81",x"CD",x"81",x"27", -- 0x0238
    x"CD",x"40",x"25",x"CD",x"00",x"1C",x"CD",x"50", -- 0x0240
    x"30",x"CD",x"A0",x"02",x"3A",x"97",x"82",x"A7", -- 0x0248
    x"C4",x"B5",x"06",x"3A",x"00",x"88",x"FD",x"E1", -- 0x0250
    x"DD",x"E1",x"C1",x"D1",x"E1",x"3E",x"01",x"32", -- 0x0258
    x"08",x"B8",x"F1",x"ED",x"45",x"3D",x"32",x"97", -- 0x0260
    x"82",x"C3",x"F0",x"01",x"21",x"5E",x"82",x"11", -- 0x0268
    x"5F",x"82",x"01",x"04",x"00",x"70",x"ED",x"B0", -- 0x0270
    x"AF",x"32",x"5C",x"82",x"CD",x"E6",x"05",x"C3", -- 0x0278
    x"53",x"02",x"3A",x"5D",x"82",x"FE",x"05",x"C2", -- 0x0280
    x"A7",x"01",x"21",x"63",x"82",x"11",x"64",x"82", -- 0x0288
    x"01",x"04",x"00",x"70",x"ED",x"B0",x"AF",x"32", -- 0x0290
    x"5D",x"82",x"CD",x"E6",x"05",x"C3",x"53",x"02", -- 0x0298
    x"2A",x"9D",x"82",x"7C",x"B5",x"C8",x"2B",x"22", -- 0x02A0
    x"9D",x"82",x"7C",x"B5",x"C0",x"32",x"AE",x"83", -- 0x02A8
    x"C9",x"AF",x"32",x"08",x"B8",x"32",x"05",x"88", -- 0x02B0
    x"32",x"10",x"B8",x"32",x"0C",x"B8",x"21",x"00", -- 0x02B8
    x"80",x"11",x"01",x"80",x"01",x"FF",x"07",x"75", -- 0x02C0
    x"ED",x"B0",x"21",x"00",x"B0",x"01",x"00",x"00", -- 0x02C8
    x"71",x"2C",x"10",x"FC",x"3A",x"02",x"E0",x"11", -- 0x02D0
    x"D6",x"0E",x"E6",x"03",x"83",x"5F",x"30",x"01", -- 0x02D8
    x"14",x"1A",x"32",x"E4",x"83",x"3A",x"04",x"E0", -- 0x02E0
    x"67",x"CB",x"5C",x"28",x"05",x"3E",x"01",x"32", -- 0x02E8
    x"C2",x"83",x"7C",x"E6",x"06",x"32",x"D4",x"83", -- 0x02F0
    x"21",x"E0",x"0E",x"11",x"EB",x"83",x"01",x"12", -- 0x02F8
    x"00",x"ED",x"B0",x"CD",x"BC",x"20",x"3E",x"01", -- 0x0300
    x"32",x"70",x"83",x"32",x"08",x"B8",x"FF",x"AF", -- 0x0308
    x"32",x"01",x"B0",x"3E",x"06",x"32",x"03",x"B0", -- 0x0310
    x"21",x"00",x"01",x"22",x"C7",x"83",x"3E",x"15", -- 0x0318
    x"32",x"81",x"83",x"21",x"87",x"0F",x"11",x"00", -- 0x0320
    x"84",x"01",x"20",x"00",x"ED",x"B0",x"21",x"06", -- 0x0328
    x"E0",x"36",x"9B",x"21",x"06",x"D0",x"36",x"88", -- 0x0330
    x"3E",x"18",x"32",x"D9",x"83",x"32",x"02",x"D0", -- 0x0338
    x"AF",x"CD",x"A7",x"07",x"3A",x"D9",x"83",x"E6", -- 0x0340
    x"EF",x"32",x"D9",x"83",x"32",x"02",x"D0",x"3E", -- 0x0348
    x"FF",x"CD",x"A7",x"07",x"3A",x"D6",x"83",x"FE", -- 0x0350
    x"02",x"D4",x"74",x"0C",x"CD",x"42",x"0B",x"3A", -- 0x0358
    x"D6",x"83",x"3D",x"C4",x"8A",x"0B",x"CD",x"98", -- 0x0360
    x"33",x"3E",x"02",x"21",x"54",x"82",x"77",x"23", -- 0x0368
    x"77",x"3E",x"09",x"23",x"77",x"23",x"77",x"23", -- 0x0370
    x"77",x"23",x"77",x"2A",x"C7",x"83",x"7C",x"B5", -- 0x0378
    x"2B",x"20",x"FB",x"3A",x"FE",x"83",x"B7",x"C2", -- 0x0380
    x"1E",x"04",x"3A",x"B3",x"83",x"B7",x"20",x"C4", -- 0x0388
    x"3A",x"02",x"E0",x"07",x"30",x"07",x"07",x"38", -- 0x0390
    x"BB",x"0E",x"02",x"18",x"02",x"0E",x"01",x"3A", -- 0x0398
    x"E1",x"83",x"B9",x"38",x"AF",x"91",x"27",x"32", -- 0x03A0
    x"E1",x"83",x"79",x"32",x"70",x"83",x"21",x"00", -- 0x03A8
    x"85",x"11",x"01",x"85",x"01",x"FF",x"01",x"75", -- 0x03B0
    x"ED",x"B0",x"32",x"FE",x"83",x"3E",x"01",x"32", -- 0x03B8
    x"FD",x"83",x"32",x"B3",x"83",x"67",x"6F",x"32", -- 0x03C0
    x"B7",x"83",x"22",x"B8",x"83",x"CD",x"2D",x"0B", -- 0x03C8
    x"3E",x"03",x"32",x"3D",x"80",x"CD",x"EC",x"07", -- 0x03D0
    x"AF",x"32",x"71",x"80",x"DF",x"3E",x"09",x"DF", -- 0x03D8
    x"3E",x"0A",x"DF",x"3E",x"0B",x"DF",x"21",x"20", -- 0x03E0
    x"00",x"22",x"9D",x"82",x"21",x"A0",x"01",x"22", -- 0x03E8
    x"82",x"83",x"21",x"00",x"00",x"22",x"D2",x"83", -- 0x03F0
    x"CD",x"F9",x"07",x"FF",x"CD",x"C6",x"32",x"AF", -- 0x03F8
    x"67",x"6F",x"32",x"2F",x"84",x"32",x"2D",x"84", -- 0x0400
    x"22",x"93",x"82",x"21",x"40",x"84",x"11",x"41", -- 0x0408
    x"84",x"01",x"4F",x"00",x"70",x"ED",x"B0",x"32", -- 0x0410
    x"04",x"80",x"3C",x"32",x"5A",x"82",x"3A",x"EA", -- 0x0418
    x"83",x"B7",x"C2",x"6A",x"04",x"3A",x"CD",x"83", -- 0x0420
    x"B7",x"20",x"0D",x"3A",x"FE",x"83",x"3D",x"28", -- 0x0428
    x"04",x"FF",x"CD",x"01",x"07",x"CD",x"42",x"0B", -- 0x0430
    x"3A",x"6D",x"82",x"A7",x"C4",x"03",x"06",x"CD", -- 0x0438
    x"65",x"09",x"32",x"EA",x"83",x"CD",x"39",x"0A", -- 0x0440
    x"21",x"9E",x"83",x"36",x"20",x"2D",x"36",x"10", -- 0x0448
    x"2D",x"36",x"20",x"3A",x"FE",x"83",x"3D",x"C4", -- 0x0450
    x"D4",x"07",x"AF",x"32",x"6D",x"82",x"3A",x"CD", -- 0x0458
    x"83",x"32",x"B6",x"83",x"CD",x"6B",x"0A",x"C3", -- 0x0460
    x"7B",x"03",x"CD",x"42",x"0B",x"3A",x"CE",x"83", -- 0x0468
    x"B7",x"CA",x"7B",x"03",x"CD",x"17",x"08",x"CD", -- 0x0470
    x"F9",x"07",x"AF",x"21",x"9A",x"83",x"77",x"2C", -- 0x0478
    x"77",x"32",x"CC",x"83",x"32",x"EA",x"83",x"21", -- 0x0480
    x"A0",x"83",x"11",x"A1",x"83",x"01",x"0D",x"00", -- 0x0488
    x"77",x"ED",x"B0",x"3E",x"80",x"DF",x"3A",x"CF", -- 0x0490
    x"83",x"B7",x"20",x"06",x"CD",x"45",x"08",x"C3", -- 0x0498
    x"7B",x"03",x"CD",x"35",x"08",x"3E",x"0C",x"DF", -- 0x04A0
    x"3E",x"0D",x"DF",x"2A",x"C5",x"83",x"2B",x"22", -- 0x04A8
    x"C5",x"83",x"7C",x"B5",x"20",x"F8",x"3A",x"FE", -- 0x04B0
    x"83",x"3D",x"CA",x"5A",x"05",x"3A",x"FD",x"83", -- 0x04B8
    x"3D",x"C2",x"06",x"05",x"21",x"C9",x"83",x"36", -- 0x04C0
    x"01",x"23",x"7E",x"B7",x"C2",x"47",x"05",x"FF", -- 0x04C8
    x"CD",x"45",x"08",x"3E",x"01",x"32",x"FE",x"83", -- 0x04D0
    x"32",x"5C",x"82",x"21",x"5E",x"82",x"11",x"5F", -- 0x04D8
    x"82",x"01",x"04",x"00",x"36",x"00",x"ED",x"B0", -- 0x04E0
    x"21",x"00",x"86",x"11",x"FF",x"80",x"01",x"B7", -- 0x04E8
    x"00",x"ED",x"B0",x"21",x"C0",x"85",x"11",x"0C", -- 0x04F0
    x"80",x"01",x"2B",x"00",x"ED",x"B0",x"3E",x"01", -- 0x04F8
    x"32",x"3F",x"80",x"C3",x"7B",x"03",x"21",x"CA", -- 0x0500
    x"83",x"36",x"01",x"2B",x"7E",x"B7",x"C2",x"6A", -- 0x0508
    x"05",x"FF",x"CD",x"45",x"08",x"3E",x"01",x"32", -- 0x0510
    x"FE",x"83",x"32",x"5D",x"82",x"21",x"63",x"82", -- 0x0518
    x"11",x"64",x"82",x"01",x"04",x"00",x"70",x"ED", -- 0x0520
    x"B0",x"21",x"C0",x"86",x"11",x"0C",x"80",x"01", -- 0x0528
    x"2B",x"00",x"ED",x"B0",x"3E",x"01",x"32",x"3F", -- 0x0530
    x"80",x"21",x"00",x"85",x"11",x"FF",x"80",x"01", -- 0x0538
    x"B7",x"00",x"ED",x"B0",x"C3",x"7B",x"03",x"AF", -- 0x0540
    x"32",x"5C",x"82",x"21",x"5E",x"82",x"11",x"5F", -- 0x0548
    x"82",x"01",x"04",x"00",x"70",x"ED",x"B0",x"C3", -- 0x0550
    x"7A",x"05",x"AF",x"32",x"5C",x"82",x"21",x"5E", -- 0x0558
    x"82",x"11",x"5F",x"82",x"01",x"04",x"00",x"70", -- 0x0560
    x"ED",x"B0",x"AF",x"32",x"5D",x"82",x"21",x"63", -- 0x0568
    x"82",x"11",x"64",x"82",x"01",x"04",x"00",x"70", -- 0x0570
    x"ED",x"B0",x"FF",x"CD",x"F9",x"07",x"CD",x"8A", -- 0x0578
    x"0B",x"CD",x"B3",x"0E",x"CD",x"42",x"0B",x"21", -- 0x0580
    x"00",x"81",x"11",x"01",x"81",x"01",x"5F",x"01", -- 0x0588
    x"75",x"ED",x"B0",x"21",x"00",x"80",x"11",x"01", -- 0x0590
    x"80",x"01",x"04",x"00",x"70",x"ED",x"B0",x"21", -- 0x0598
    x"0C",x"80",x"11",x"0D",x"80",x"01",x"2E",x"00", -- 0x05A0
    x"70",x"ED",x"B0",x"AF",x"32",x"C3",x"83",x"32", -- 0x05A8
    x"FE",x"83",x"32",x"BF",x"83",x"21",x"C9",x"83", -- 0x05B0
    x"77",x"2C",x"77",x"67",x"6F",x"32",x"10",x"B8", -- 0x05B8
    x"32",x"0C",x"B8",x"22",x"93",x"82",x"32",x"BB", -- 0x05C0
    x"83",x"32",x"CB",x"83",x"32",x"D8",x"83",x"32", -- 0x05C8
    x"C4",x"83",x"32",x"BA",x"83",x"32",x"95",x"82", -- 0x05D0
    x"32",x"5B",x"82",x"3E",x"03",x"32",x"D6",x"83", -- 0x05D8
    x"CD",x"FE",x"07",x"C3",x"7B",x"03",x"3E",x"01", -- 0x05E0
    x"32",x"6D",x"82",x"32",x"5A",x"82",x"32",x"CD", -- 0x05E8
    x"83",x"AF",x"32",x"5B",x"82",x"32",x"EA",x"83", -- 0x05F0
    x"3E",x"FF",x"32",x"97",x"82",x"3E",x"40",x"32", -- 0x05F8
    x"98",x"82",x"C9",x"3E",x"10",x"DF",x"3E",x"30", -- 0x0600
    x"DF",x"3A",x"FD",x"83",x"3D",x"20",x"0C",x"21", -- 0x0608
    x"93",x"82",x"34",x"7E",x"D6",x"05",x"20",x"0D", -- 0x0610
    x"77",x"18",x"0A",x"21",x"94",x"82",x"34",x"7E", -- 0x0618
    x"D6",x"05",x"20",x"01",x"77",x"CD",x"3C",x"06", -- 0x0620
    x"CD",x"5E",x"06",x"CD",x"C6",x"32",x"CD",x"8B", -- 0x0628
    x"2A",x"3E",x"01",x"32",x"80",x"83",x"11",x"00", -- 0x0630
    x"01",x"C3",x"03",x"09",x"CD",x"F9",x"07",x"21", -- 0x0638
    x"9A",x"83",x"AF",x"77",x"2C",x"77",x"3C",x"32", -- 0x0640
    x"CC",x"83",x"3E",x"20",x"21",x"06",x"A8",x"CD", -- 0x0648
    x"8C",x"07",x"2C",x"2C",x"CD",x"8C",x"07",x"0E", -- 0x0650
    x"0A",x"09",x"3D",x"20",x"F2",x"C9",x"21",x"0C", -- 0x0658
    x"80",x"11",x"0D",x"80",x"01",x"2B",x"00",x"70", -- 0x0660
    x"ED",x"B0",x"21",x"0C",x"80",x"11",x"0C",x"B0", -- 0x0668
    x"01",x"2B",x"00",x"ED",x"B0",x"21",x"00",x"81", -- 0x0670
    x"11",x"01",x"81",x"01",x"62",x"00",x"36",x"00", -- 0x0678
    x"ED",x"B0",x"C9",x"21",x"64",x"AB",x"CD",x"A8", -- 0x0680
    x"06",x"21",x"A4",x"AA",x"CD",x"A8",x"06",x"21", -- 0x0688
    x"E4",x"A9",x"CD",x"A8",x"06",x"21",x"24",x"A9", -- 0x0690
    x"CD",x"A8",x"06",x"21",x"64",x"A8",x"CD",x"A8", -- 0x0698
    x"06",x"AF",x"32",x"2F",x"84",x"C3",x"82",x"0A", -- 0x06A0
    x"3E",x"10",x"77",x"23",x"77",x"01",x"1F",x"00", -- 0x06A8
    x"09",x"77",x"23",x"77",x"C9",x"FE",x"C0",x"CA", -- 0x06B0
    x"D4",x"06",x"FE",x"90",x"CA",x"DA",x"06",x"FE", -- 0x06B8
    x"70",x"CA",x"E0",x"06",x"FE",x"50",x"CA",x"E6", -- 0x06C0
    x"06",x"FE",x"30",x"CA",x"EC",x"06",x"FE",x"10", -- 0x06C8
    x"CA",x"83",x"06",x"C9",x"21",x"64",x"AB",x"C3", -- 0x06D0
    x"F2",x"06",x"21",x"A4",x"AA",x"C3",x"F2",x"06", -- 0x06D8
    x"21",x"E4",x"A9",x"C3",x"F2",x"06",x"21",x"24", -- 0x06E0
    x"A9",x"C3",x"F2",x"06",x"21",x"64",x"A8",x"C3", -- 0x06E8
    x"F2",x"06",x"36",x"FC",x"23",x"36",x"FD",x"01", -- 0x06F0
    x"1F",x"00",x"09",x"36",x"FE",x"23",x"36",x"FF", -- 0x06F8
    x"C9",x"3A",x"FD",x"83",x"3D",x"20",x"32",x"21", -- 0x0700
    x"0C",x"80",x"11",x"C0",x"85",x"01",x"2B",x"00", -- 0x0708
    x"ED",x"B0",x"21",x"FF",x"80",x"11",x"00",x"86", -- 0x0710
    x"01",x"B7",x"00",x"ED",x"B0",x"21",x"C0",x"86", -- 0x0718
    x"11",x"0C",x"80",x"01",x"2B",x"00",x"ED",x"B0", -- 0x0720
    x"3E",x"01",x"32",x"3F",x"80",x"21",x"00",x"85", -- 0x0728
    x"11",x"FF",x"80",x"01",x"B7",x"00",x"ED",x"B0", -- 0x0730
    x"C9",x"21",x"FF",x"80",x"11",x"00",x"85",x"01", -- 0x0738
    x"B7",x"00",x"ED",x"B0",x"21",x"0C",x"80",x"11", -- 0x0740
    x"C0",x"86",x"01",x"2B",x"00",x"ED",x"B0",x"21", -- 0x0748
    x"00",x"86",x"11",x"FF",x"80",x"01",x"B7",x"00", -- 0x0750
    x"ED",x"B0",x"21",x"C0",x"85",x"11",x"0C",x"80", -- 0x0758
    x"01",x"2B",x"00",x"ED",x"B0",x"3E",x"01",x"32", -- 0x0760
    x"3F",x"80",x"3A",x"95",x"82",x"A7",x"C0",x"AF", -- 0x0768
    x"32",x"5B",x"82",x"3E",x"01",x"32",x"95",x"82", -- 0x0770
    x"C9",x"21",x"02",x"A8",x"11",x"10",x"20",x"0E", -- 0x0778
    x"04",x"06",x"1C",x"73",x"23",x"10",x"FC",x"09", -- 0x0780
    x"15",x"20",x"F6",x"C9",x"01",x"10",x"0A",x"71", -- 0x0788
    x"23",x"10",x"FC",x"C9",x"21",x"08",x"A8",x"11", -- 0x0790
    x"10",x"20",x"0E",x"0A",x"06",x"16",x"73",x"23", -- 0x0798
    x"10",x"FC",x"09",x"15",x"20",x"F6",x"C9",x"32", -- 0x07A0
    x"00",x"D0",x"3A",x"D9",x"83",x"E6",x"F7",x"32", -- 0x07A8
    x"02",x"D0",x"00",x"00",x"00",x"00",x"3A",x"D9", -- 0x07B0
    x"83",x"F6",x"08",x"32",x"02",x"D0",x"C9",x"21", -- 0x07B8
    x"00",x"83",x"7E",x"B7",x"C8",x"35",x"4F",x"2C", -- 0x07C0
    x"7E",x"CD",x"A7",x"07",x"54",x"5D",x"2C",x"06", -- 0x07C8
    x"00",x"ED",x"B0",x"C9",x"3A",x"FD",x"83",x"3D", -- 0x07D0
    x"CA",x"E1",x"07",x"3E",x"01",x"32",x"5B",x"82", -- 0x07D8
    x"C9",x"3A",x"6D",x"82",x"A7",x"C8",x"3E",x"01", -- 0x07E0
    x"32",x"5B",x"82",x"C9",x"21",x"00",x"83",x"11", -- 0x07E8
    x"01",x"83",x"01",x"2F",x"00",x"70",x"ED",x"B0", -- 0x07F0
    x"C9",x"3A",x"FE",x"83",x"3D",x"C8",x"AF",x"21", -- 0x07F8
    x"44",x"80",x"11",x"45",x"80",x"01",x"1F",x"00", -- 0x0800
    x"70",x"ED",x"B0",x"21",x"20",x"84",x"11",x"21", -- 0x0808
    x"84",x"0E",x"0B",x"77",x"ED",x"B0",x"C9",x"21", -- 0x0810
    x"44",x"80",x"AF",x"36",x"01",x"2C",x"77",x"2C", -- 0x0818
    x"2C",x"77",x"3A",x"FE",x"83",x"FE",x"02",x"C0", -- 0x0820
    x"21",x"40",x"00",x"22",x"D2",x"83",x"21",x"40", -- 0x0828
    x"00",x"22",x"DA",x"83",x"C9",x"21",x"50",x"A8", -- 0x0830
    x"CD",x"6B",x"2A",x"21",x"70",x"AA",x"11",x"D6", -- 0x0838
    x"0F",x"06",x"09",x"EF",x"C9",x"AF",x"32",x"71", -- 0x0840
    x"83",x"3A",x"FE",x"83",x"3D",x"C8",x"3A",x"FD", -- 0x0848
    x"83",x"EE",x"03",x"32",x"FD",x"83",x"21",x"B8", -- 0x0850
    x"83",x"3D",x"28",x"01",x"2C",x"7E",x"32",x"B7", -- 0x0858
    x"83",x"AF",x"32",x"B6",x"83",x"3C",x"32",x"5A", -- 0x0860
    x"82",x"3A",x"C2",x"83",x"B7",x"C8",x"3A",x"CB", -- 0x0868
    x"83",x"EE",x"01",x"32",x"CB",x"83",x"67",x"32", -- 0x0870
    x"10",x"B8",x"32",x"0C",x"B8",x"C9",x"21",x"51", -- 0x0878
    x"AA",x"11",x"04",x"10",x"06",x"04",x"EF",x"11", -- 0x0880
    x"DA",x"0F",x"06",x"05",x"EF",x"3E",x"01",x"32", -- 0x0888
    x"04",x"80",x"C9",x"3A",x"CD",x"83",x"B7",x"C0", -- 0x0890
    x"3A",x"04",x"80",x"B7",x"C0",x"3A",x"AE",x"83", -- 0x0898
    x"B7",x"20",x"07",x"3C",x"32",x"AE",x"83",x"3E", -- 0x08A0
    x"06",x"DF",x"CD",x"DD",x"0A",x"3A",x"DF",x"83", -- 0x08A8
    x"B7",x"20",x"35",x"21",x"DC",x"83",x"35",x"C0", -- 0x08B0
    x"36",x"20",x"23",x"7E",x"B7",x"CA",x"7E",x"08", -- 0x08B8
    x"3D",x"77",x"2C",x"7E",x"3D",x"27",x"77",x"2D", -- 0x08C0
    x"FE",x"10",x"20",x"07",x"3E",x"05",x"DF",x"AF", -- 0x08C8
    x"32",x"3F",x"80",x"66",x"7C",x"E6",x"03",x"4F", -- 0x08D0
    x"AC",x"07",x"07",x"6F",x"26",x"00",x"29",x"11", -- 0x08D8
    x"DF",x"A8",x"19",x"3E",x"10",x"91",x"77",x"C9", -- 0x08E0
    x"3A",x"E0",x"83",x"B7",x"C0",x"3C",x"32",x"E0", -- 0x08E8
    x"83",x"21",x"51",x"AA",x"11",x"04",x"10",x"06", -- 0x08F0
    x"05",x"EF",x"3A",x"DE",x"83",x"5F",x"16",x"00", -- 0x08F8
    x"CD",x"C3",x"0B",x"3A",x"FE",x"83",x"B7",x"C8", -- 0x0900
    x"3A",x"FD",x"83",x"3D",x"28",x"05",x"21",x"EB", -- 0x0908
    x"83",x"18",x"03",x"21",x"ED",x"83",x"7B",x"86", -- 0x0910
    x"27",x"77",x"5F",x"23",x"7A",x"8E",x"27",x"77", -- 0x0918
    x"57",x"3A",x"FD",x"83",x"3D",x"20",x"09",x"01", -- 0x0920
    x"E7",x"83",x"0A",x"B7",x"20",x"2B",x"18",x"07", -- 0x0928
    x"01",x"E8",x"83",x"0A",x"B7",x"20",x"22",x"2A", -- 0x0930
    x"DE",x"0E",x"ED",x"52",x"28",x"02",x"30",x"19", -- 0x0938
    x"32",x"CF",x"83",x"3C",x"02",x"0D",x"0D",x"0A", -- 0x0940
    x"3C",x"02",x"21",x"DE",x"AB",x"01",x"E0",x"FF", -- 0x0948
    x"09",x"3D",x"20",x"FC",x"36",x"4D",x"3E",x"07", -- 0x0950
    x"DF",x"2A",x"EF",x"83",x"B7",x"ED",x"52",x"D0", -- 0x0958
    x"ED",x"53",x"EF",x"83",x"C9",x"AF",x"32",x"CE", -- 0x0960
    x"83",x"3A",x"CD",x"83",x"B7",x"20",x"04",x"AF", -- 0x0968
    x"32",x"CF",x"83",x"3A",x"FE",x"83",x"B7",x"28", -- 0x0970
    x"74",x"3A",x"FD",x"83",x"3D",x"20",x"05",x"21", -- 0x0978
    x"E5",x"83",x"18",x"03",x"21",x"E6",x"83",x"3A", -- 0x0980
    x"CD",x"83",x"B7",x"20",x"08",x"35",x"20",x"05", -- 0x0988
    x"3E",x"01",x"32",x"CF",x"83",x"CD",x"DB",x"29", -- 0x0990
    x"3A",x"CD",x"83",x"B7",x"20",x"0A",x"3C",x"32", -- 0x0998
    x"B5",x"83",x"21",x"50",x"A8",x"CD",x"6B",x"2A", -- 0x09A0
    x"3A",x"6C",x"82",x"EE",x"01",x"32",x"B5",x"83", -- 0x09A8
    x"3A",x"FD",x"83",x"3D",x"C2",x"F5",x"09",x"21", -- 0x09B0
    x"5E",x"82",x"CD",x"FE",x"09",x"3A",x"5A",x"82", -- 0x09B8
    x"A7",x"28",x"0A",x"CD",x"C6",x"32",x"CD",x"23", -- 0x09C0
    x"20",x"AF",x"32",x"5A",x"82",x"21",x"44",x"80", -- 0x09C8
    x"36",x"80",x"2C",x"36",x"1E",x"2C",x"36",x"03", -- 0x09D0
    x"2C",x"36",x"E0",x"AF",x"32",x"CD",x"83",x"32", -- 0x09D8
    x"2D",x"84",x"32",x"2C",x"84",x"32",x"69",x"82", -- 0x09E0
    x"3C",x"32",x"C3",x"83",x"C9",x"3A",x"CD",x"83", -- 0x09E8
    x"B7",x"C8",x"C3",x"CD",x"09",x"21",x"63",x"82", -- 0x09F0
    x"CD",x"FE",x"09",x"C3",x"BD",x"09",x"AF",x"B6", -- 0x09F8
    x"11",x"64",x"AB",x"C4",x"28",x"0A",x"23",x"AF", -- 0x0A00
    x"B6",x"11",x"A4",x"AA",x"C4",x"28",x"0A",x"23", -- 0x0A08
    x"AF",x"B6",x"11",x"E4",x"A9",x"C4",x"28",x"0A", -- 0x0A10
    x"23",x"AF",x"B6",x"11",x"24",x"A9",x"C4",x"28", -- 0x0A18
    x"0A",x"23",x"AF",x"B6",x"11",x"64",x"A8",x"C8", -- 0x0A20
    x"EB",x"36",x"6C",x"23",x"36",x"6D",x"01",x"1F", -- 0x0A28
    x"00",x"09",x"36",x"6E",x"23",x"36",x"6F",x"EB", -- 0x0A30
    x"C9",x"3A",x"E4",x"83",x"3C",x"C8",x"3A",x"FE", -- 0x0A38
    x"83",x"B7",x"20",x"05",x"21",x"E4",x"83",x"18", -- 0x0A40
    x"0E",x"3A",x"FD",x"83",x"3D",x"20",x"05",x"21", -- 0x0A48
    x"E5",x"83",x"18",x"03",x"21",x"E6",x"83",x"46", -- 0x0A50
    x"78",x"B7",x"3E",x"4D",x"11",x"E0",x"FF",x"21", -- 0x0A58
    x"BE",x"AB",x"28",x"04",x"77",x"19",x"10",x"FC", -- 0x0A60
    x"36",x"10",x"C9",x"3A",x"B7",x"83",x"21",x"7E", -- 0x0A68
    x"A8",x"11",x"20",x"00",x"FE",x"0F",x"38",x"02", -- 0x0A70
    x"3E",x"0F",x"47",x"0E",x"4C",x"71",x"19",x"10", -- 0x0A78
    x"FC",x"C9",x"AF",x"32",x"CC",x"83",x"21",x"B8", -- 0x0A80
    x"83",x"3A",x"FD",x"83",x"3D",x"28",x"01",x"2C", -- 0x0A88
    x"34",x"7E",x"32",x"B7",x"83",x"FE",x"10",x"D0", -- 0x0A90
    x"26",x"00",x"11",x"5E",x"A8",x"87",x"87",x"87", -- 0x0A98
    x"87",x"6F",x"29",x"19",x"36",x"4C",x"C9",x"06", -- 0x0AA0
    x"05",x"21",x"F2",x"83",x"7A",x"BE",x"38",x"27", -- 0x0AA8
    x"28",x"19",x"78",x"3D",x"28",x"0F",x"87",x"4F", -- 0x0AB0
    x"06",x"00",x"D5",x"11",x"FA",x"83",x"21",x"F8", -- 0x0AB8
    x"83",x"ED",x"B8",x"EB",x"D1",x"72",x"2D",x"73", -- 0x0AC0
    x"87",x"3C",x"C9",x"2D",x"7E",x"2C",x"BB",x"38", -- 0x0AC8
    x"E1",x"20",x"04",x"78",x"3D",x"28",x"F1",x"2C", -- 0x0AD0
    x"2C",x"10",x"D1",x"AF",x"C9",x"3A",x"2D",x"84", -- 0x0AD8
    x"B7",x"C0",x"3C",x"32",x"2D",x"84",x"3E",x"03", -- 0x0AE0
    x"32",x"3F",x"80",x"AF",x"32",x"E0",x"83",x"21", -- 0x0AE8
    x"BF",x"A8",x"11",x"04",x"10",x"06",x"04",x"EF", -- 0x0AF0
    x"21",x"DF",x"A8",x"11",x"20",x"00",x"01",x"0C", -- 0x0AF8
    x"0F",x"71",x"19",x"10",x"FC",x"21",x"20",x"3C", -- 0x0B00
    x"22",x"DC",x"83",x"3E",x"60",x"32",x"DE",x"83", -- 0x0B08
    x"C9",x"E5",x"D5",x"21",x"00",x"84",x"35",x"20", -- 0x0B10
    x"02",x"36",x"1F",x"54",x"5E",x"7B",x"C6",x"0D", -- 0x0B18
    x"FE",x"20",x"38",x"02",x"D6",x"1F",x"6F",x"1A", -- 0x0B20
    x"AE",x"77",x"D1",x"E1",x"C9",x"21",x"00",x"00", -- 0x0B28
    x"22",x"ED",x"83",x"22",x"EB",x"83",x"22",x"E7", -- 0x0B30
    x"83",x"3A",x"E4",x"83",x"67",x"6F",x"22",x"E5", -- 0x0B38
    x"83",x"C9",x"11",x"AA",x"0F",x"21",x"60",x"AA", -- 0x0B40
    x"06",x"08",x"EF",x"21",x"41",x"AA",x"ED",x"5B", -- 0x0B48
    x"EF",x"83",x"CD",x"B8",x"0B",x"3E",x"01",x"21", -- 0x0B50
    x"20",x"AB",x"CD",x"CC",x"0B",x"11",x"A7",x"0F", -- 0x0B58
    x"06",x"03",x"EF",x"21",x"41",x"AB",x"ED",x"5B", -- 0x0B60
    x"ED",x"83",x"CD",x"B8",x"0B",x"3A",x"70",x"83", -- 0x0B68
    x"3D",x"C8",x"3E",x"02",x"21",x"00",x"A9",x"CD", -- 0x0B70
    x"CC",x"0B",x"11",x"A7",x"0F",x"06",x"03",x"EF", -- 0x0B78
    x"21",x"21",x"A9",x"ED",x"5B",x"EB",x"83",x"C3", -- 0x0B80
    x"B8",x"0B",x"3A",x"B4",x"83",x"B7",x"20",x"11", -- 0x0B88
    x"3C",x"32",x"B4",x"83",x"21",x"1F",x"A8",x"11", -- 0x0B90
    x"20",x"00",x"01",x"10",x"20",x"71",x"19",x"10", -- 0x0B98
    x"FC",x"11",x"FE",x"0F",x"21",x"7F",x"A9",x"06", -- 0x0BA0
    x"06",x"EF",x"3E",x"01",x"32",x"3F",x"80",x"21", -- 0x0BA8
    x"9F",x"A8",x"3A",x"E1",x"83",x"C3",x"C3",x"0B", -- 0x0BB0
    x"CD",x"BE",x"0B",x"AF",x"18",x"0E",x"7A",x"CD", -- 0x0BB8
    x"C3",x"0B",x"7B",x"4F",x"0F",x"0F",x"0F",x"0F", -- 0x0BC0
    x"CD",x"CC",x"0B",x"79",x"E6",x"0F",x"77",x"7D", -- 0x0BC8
    x"D6",x"20",x"6F",x"D0",x"25",x"C9",x"21",x"D8", -- 0x0BD0
    x"83",x"35",x"2D",x"AF",x"77",x"32",x"B3",x"83", -- 0x0BD8
    x"CD",x"79",x"07",x"3E",x"03",x"32",x"19",x"80", -- 0x0BE0
    x"21",x"1F",x"80",x"06",x"05",x"AF",x"77",x"2C", -- 0x0BE8
    x"2C",x"2C",x"2C",x"10",x"F9",x"CD",x"60",x"0C", -- 0x0BF0
    x"21",x"AC",x"AA",x"11",x"AD",x"0F",x"06",x"0D", -- 0x0BF8
    x"EF",x"3E",x"01",x"26",x"AA",x"ED",x"47",x"87", -- 0x0C00
    x"C6",x"CD",x"6F",x"ED",x"57",x"CD",x"CC",x"0B", -- 0x0C08
    x"ED",x"57",x"08",x"06",x"03",x"EF",x"D9",x"21", -- 0x0C10
    x"EF",x"83",x"08",x"47",x"2C",x"2C",x"10",x"FC", -- 0x0C18
    x"5E",x"2C",x"56",x"26",x"A9",x"87",x"C6",x"ED", -- 0x0C20
    x"6F",x"CD",x"B8",x"0B",x"11",x"4B",x"10",x"06", -- 0x0C28
    x"04",x"EF",x"ED",x"57",x"D9",x"3C",x"FE",x"06", -- 0x0C30
    x"20",x"C9",x"11",x"DF",x"0F",x"21",x"3C",x"AB", -- 0x0C38
    x"06",x"13",x"AF",x"32",x"39",x"80",x"EF",x"C9", -- 0x0C40
    x"7A",x"CD",x"4D",x"0C",x"7B",x"4F",x"E6",x"0F", -- 0x0C48
    x"CD",x"58",x"0C",x"79",x"0F",x"0F",x"0F",x"0F", -- 0x0C50
    x"77",x"7D",x"D6",x"20",x"6F",x"D0",x"25",x"C9", -- 0x0C58
    x"26",x"80",x"ED",x"4B",x"FB",x"83",x"11",x"04", -- 0x0C60
    x"30",x"CD",x"6D",x"0C",x"48",x"7A",x"91",x"BA", -- 0x0C68
    x"C8",x"6F",x"73",x"C9",x"3A",x"D8",x"83",x"B7", -- 0x0C70
    x"C0",x"3A",x"D6",x"83",x"FE",x"03",x"CA",x"D6", -- 0x0C78
    x"0B",x"3A",x"E1",x"83",x"B7",x"C2",x"A6",x"0C", -- 0x0C80
    x"3A",x"D6",x"83",x"FE",x"04",x"CA",x"00",x"18", -- 0x0C88
    x"FE",x"02",x"CA",x"9B",x"3E",x"FE",x"05",x"C0", -- 0x0C90
    x"21",x"D8",x"83",x"36",x"30",x"2D",x"AF",x"77", -- 0x0C98
    x"32",x"15",x"80",x"C3",x"3A",x"0C",x"CD",x"F9", -- 0x0CA0
    x"07",x"3A",x"BA",x"83",x"B7",x"C0",x"67",x"6F", -- 0x0CA8
    x"22",x"93",x"82",x"22",x"B3",x"81",x"32",x"5B", -- 0x0CB0
    x"82",x"32",x"9A",x"82",x"3C",x"32",x"BA",x"83", -- 0x0CB8
    x"CD",x"C6",x"32",x"CD",x"17",x"08",x"CD",x"79", -- 0x0CC0
    x"07",x"CD",x"5E",x"06",x"3E",x"04",x"32",x"1B", -- 0x0CC8
    x"80",x"3E",x"06",x"32",x"29",x"80",x"21",x"28", -- 0x0CD0
    x"AA",x"11",x"0D",x"10",x"06",x"04",x"EF",x"21", -- 0x0CD8
    x"AD",x"AA",x"13",x"06",x"0C",x"EF",x"CD",x"13", -- 0x0CE0
    x"0D",x"21",x"74",x"AB",x"11",x"1E",x"10",x"06", -- 0x0CE8
    x"03",x"EF",x"11",x"39",x"10",x"06",x"06",x"EF", -- 0x0CF0
    x"11",x"3F",x"10",x"06",x"05",x"EF",x"13",x"06", -- 0x0CF8
    x"07",x"EF",x"21",x"94",x"A9",x"ED",x"5B",x"DE", -- 0x0D00
    x"0E",x"CD",x"B8",x"0B",x"11",x"4B",x"10",x"06", -- 0x0D08
    x"04",x"EF",x"C9",x"3A",x"E1",x"83",x"11",x"1E", -- 0x0D10
    x"10",x"3D",x"28",x"11",x"3E",x"03",x"32",x"23", -- 0x0D18
    x"80",x"21",x"11",x"AB",x"06",x"04",x"EF",x"06", -- 0x0D20
    x"0D",x"EF",x"36",x"23",x"C9",x"21",x"F1",x"AA", -- 0x0D28
    x"06",x"04",x"EF",x"11",x"29",x"10",x"06",x"0B", -- 0x0D30
    x"EF",x"C9",x"3E",x"03",x"32",x"0D",x"80",x"32", -- 0x0D38
    x"0F",x"80",x"3A",x"BC",x"83",x"3D",x"32",x"BC", -- 0x0D40
    x"83",x"C0",x"3E",x"20",x"32",x"BC",x"83",x"3A", -- 0x0D48
    x"D7",x"83",x"87",x"16",x"00",x"5F",x"21",x"59", -- 0x0D50
    x"0D",x"19",x"E9",x"18",x"46",x"18",x"3A",x"18", -- 0x0D58
    x"2E",x"18",x"22",x"18",x"16",x"18",x"0A",x"21", -- 0x0D60
    x"06",x"AB",x"11",x"40",x"80",x"3E",x"D4",x"18", -- 0x0D68
    x"3A",x"21",x"A6",x"AA",x"11",x"44",x"80",x"3E", -- 0x0D70
    x"D8",x"18",x"30",x"21",x"46",x"AA",x"11",x"48", -- 0x0D78
    x"80",x"3E",x"DC",x"18",x"26",x"21",x"E6",x"A9", -- 0x0D80
    x"11",x"4C",x"80",x"3E",x"F4",x"18",x"1C",x"21", -- 0x0D88
    x"86",x"A9",x"11",x"50",x"80",x"3E",x"F4",x"18", -- 0x0D90
    x"12",x"21",x"26",x"A9",x"11",x"54",x"80",x"3E", -- 0x0D98
    x"F8",x"18",x"08",x"21",x"C6",x"A8",x"11",x"58", -- 0x0DA0
    x"80",x"3E",x"D8",x"01",x"1F",x"00",x"77",x"3C", -- 0x0DA8
    x"2C",x"77",x"3C",x"09",x"77",x"3C",x"2C",x"77", -- 0x0DB0
    x"EB",x"01",x"00",x"04",x"71",x"2C",x"10",x"FC", -- 0x0DB8
    x"21",x"D7",x"83",x"35",x"C0",x"36",x"07",x"AF", -- 0x0DC0
    x"32",x"BF",x"83",x"32",x"BB",x"83",x"3E",x"05", -- 0x0DC8
    x"32",x"D6",x"83",x"C9",x"3A",x"E1",x"83",x"B7", -- 0x0DD0
    x"20",x"F4",x"21",x"BF",x"83",x"7E",x"B7",x"20", -- 0x0DD8
    x"2D",x"CD",x"79",x"07",x"CD",x"5E",x"06",x"21", -- 0x0DE0
    x"40",x"80",x"01",x"03",x"07",x"11",x"00",x"81", -- 0x0DE8
    x"73",x"2C",x"2C",x"71",x"2C",x"72",x"2C",x"10", -- 0x0DF0
    x"F7",x"21",x"04",x"05",x"22",x"BD",x"83",x"21", -- 0x0DF8
    x"D7",x"83",x"36",x"07",x"21",x"BC",x"83",x"36", -- 0x0E00
    x"20",x"21",x"BF",x"83",x"34",x"C9",x"3D",x"20", -- 0x0E08
    x"5F",x"3A",x"D7",x"83",x"87",x"16",x"00",x"5F", -- 0x0E10
    x"21",x"1B",x"0E",x"19",x"E9",x"18",x"34",x"18", -- 0x0E18
    x"2B",x"18",x"22",x"18",x"19",x"18",x"10",x"18", -- 0x0E20
    x"07",x"21",x"40",x"80",x"06",x"31",x"18",x"28", -- 0x0E28
    x"21",x"44",x"80",x"06",x"49",x"18",x"21",x"21", -- 0x0E30
    x"48",x"80",x"06",x"61",x"18",x"1A",x"21",x"4C", -- 0x0E38
    x"80",x"06",x"79",x"18",x"13",x"21",x"50",x"80", -- 0x0E40
    x"06",x"91",x"18",x"0C",x"21",x"54",x"80",x"06", -- 0x0E48
    x"A9",x"18",x"05",x"21",x"58",x"80",x"06",x"C1", -- 0x0E50
    x"CD",x"98",x"0E",x"4F",x"35",x"35",x"35",x"35", -- 0x0E58
    x"7E",x"2C",x"71",x"B8",x"D0",x"36",x"1E",x"21", -- 0x0E60
    x"D7",x"83",x"35",x"C0",x"36",x"14",x"18",x"99", -- 0x0E68
    x"3D",x"C2",x"3A",x"0D",x"CD",x"98",x"0E",x"D6", -- 0x0E70
    x"03",x"4F",x"3A",x"D7",x"83",x"B7",x"CA",x"FF", -- 0x0E78
    x"0D",x"06",x"07",x"11",x"06",x"00",x"21",x"43", -- 0x0E80
    x"80",x"35",x"35",x"35",x"35",x"2D",x"2D",x"71", -- 0x0E88
    x"19",x"10",x"F6",x"3D",x"32",x"D7",x"83",x"C9", -- 0x0E90
    x"E5",x"21",x"BD",x"83",x"35",x"20",x"11",x"36", -- 0x0E98
    x"08",x"2C",x"35",x"20",x"02",x"36",x"04",x"7E", -- 0x0EA0
    x"21",x"F1",x"0E",x"85",x"6F",x"7E",x"E1",x"C9", -- 0x0EA8
    x"F1",x"F1",x"C9",x"ED",x"5B",x"ED",x"83",x"2A", -- 0x0EB0
    x"EB",x"83",x"44",x"4D",x"B7",x"ED",x"52",x"38", -- 0x0EB8
    x"05",x"D5",x"C5",x"D1",x"18",x"01",x"C5",x"CD", -- 0x0EC0
    x"A7",x"0A",x"D1",x"F5",x"CD",x"A7",x"0A",x"67", -- 0x0EC8
    x"F1",x"6F",x"22",x"FB",x"83",x"C9",x"03",x"05", -- 0x0ED0
    x"07",x"FF",x"00",x"02",x"04",x"06",x"00",x"20", -- 0x0ED8
    x"00",x"00",x"58",x"01",x"63",x"04",x"63",x"04", -- 0x0EE0
    x"05",x"02",x"97",x"01",x"58",x"01",x"27",x"01", -- 0x0EE8
    x"05",x"00",x"1F",x"20",x"21",x"20",x"25",x"26", -- 0x0EF0
    x"27",x"26",x"2C",x"2D",x"2E",x"2D",x"2F",x"30", -- 0x0EF8
    x"31",x"30",x"2C",x"2E",x"30",x"2E",x"2D",x"2F", -- 0x0F00
    x"31",x"2F",x"25",x"26",x"27",x"2C",x"2D",x"2E", -- 0x0F08
    x"2F",x"30",x"31",x"2C",x"2E",x"30",x"2D",x"2F", -- 0x0F10
    x"31",x"04",x"04",x"04",x"08",x"08",x"08",x"08", -- 0x0F18
    x"08",x"08",x"10",x"10",x"10",x"02",x"03",x"03", -- 0x0F20
    x"05",x"05",x"06",x"08",x"09",x"54",x"58",x"5A", -- 0x0F28
    x"5E",x"56",x"5C",x"03",x"03",x"06",x"08",x"10", -- 0x0F30
    x"18",x"30",x"50",x"60",x"80",x"C0",x"E0",x"05", -- 0x0F38
    x"02",x"02",x"02",x"08",x"08",x"05",x"08",x"02", -- 0x0F40
    x"08",x"08",x"08",x"0E",x"08",x"08",x"0E",x"08", -- 0x0F48
    x"0E",x"08",x"0E",x"08",x"0E",x"08",x"05",x"05", -- 0x0F50
    x"08",x"05",x"02",x"0B",x"05",x"08",x"FF",x"C0", -- 0x0F58
    x"02",x"00",x"03",x"00",x"03",x"80",x"01",x"80", -- 0x0F60
    x"02",x"80",x"02",x"00",x"02",x"00",x"02",x"80", -- 0x0F68
    x"03",x"E0",x"02",x"20",x"02",x"20",x"02",x"20", -- 0x0F70
    x"02",x"00",x"03",x"80",x"02",x"C0",x"02",x"C0", -- 0x0F78
    x"02",x"80",x"03",x"20",x"02",x"20",x"02",x"10", -- 0x0F80
    x"3B",x"8C",x"D9",x"AF",x"7F",x"3C",x"30",x"70", -- 0x0F88
    x"A9",x"47",x"E7",x"A7",x"FF",x"BC",x"36",x"10", -- 0x0F90
    x"F9",x"40",x"D2",x"D7",x"C4",x"37",x"A6",x"9B", -- 0x0F98
    x"A1",x"00",x"C7",x"AC",x"8D",x"C5",x"06",x"2B", -- 0x0FA0
    x"25",x"20",x"18",x"19",x"2B",x"23",x"13",x"1F", -- 0x0FA8
    x"22",x"15",x"10",x"22",x"11",x"1E",x"1B",x"19", -- 0x0FB0
    x"1E",x"17",x"10",x"23",x"24",x"10",x"1E",x"14", -- 0x0FB8
    x"10",x"22",x"14",x"10",x"24",x"18",x"10",x"24", -- 0x0FC0
    x"18",x"2B",x"20",x"1F",x"19",x"1E",x"24",x"10", -- 0x0FC8
    x"24",x"11",x"12",x"1C",x"15",x"2B",x"17",x"11", -- 0x0FD0
    x"1D",x"15",x"10",x"1F",x"26",x"15",x"22",x"10", -- 0x0FD8
    x"10",x"10",x"23",x"15",x"17",x"11",x"10",x"10", -- 0x0FE0
    x"4E",x"10",x"10",x"01",x"09",x"08",x"01",x"10", -- 0x0FE8
    x"10",x"10",x"19",x"1E",x"23",x"15",x"22",x"24", -- 0x0FF0
    x"10",x"13",x"1F",x"19",x"1E",x"23",x"13",x"22"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
